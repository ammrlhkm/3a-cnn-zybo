--------------------------------------------------------------------------------
-- VHDL ROM with NORMALIZED image pixels (fixed-point format)
-- Generated from: 3_tabby_cat_s_001397.ppm
-- Generated on: 2025-12-11 22:11:27
-- 
-- Image size: 24x24 RGB
-- Memory depth: 1728 values
-- Address bits: 11
--
-- Normalization applied (matches cnn_ref.py):
--   mean = 167.3929
--   std_dev = 35.3794
--   normalized = (pixel - mean) / std_dev
--
-- Fixed-point format: Q5.5 (signed)
--   Total bits: 10
--   Integer bits: 5 (including sign)
--   Fractional bits: 5
--   Range: [-16.0000, 15.9688]
--   Resolution: 0.031250
--
-- Memory layout: Interleaved RGB
--   addr = (h * 24 + w) * 3 + channel
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity input_image_rom is
    generic (
        CELL_COUNT : integer := 1728;
        ADDR_WIDTH : integer := 11;
        DATA_WIDTH : integer := 10
    );
    port (
        clk     : in  std_logic;
        addr    : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        dout    : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end entity input_image_rom;

architecture rtl of input_image_rom is
    
    type mem_type is array (0 to CELL_COUNT-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

    -- Output register for better timing (addresses SYNTH-6 warning)
    signal dout_reg : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');

    -- Normalized fixed-point pixel values
    constant mem : mem_type := (
        0 => "1110101010",  -- -2.6963
        1 => "1110011011",  -- -3.1485
        2 => "1110010111",  -- -3.2899
        3 => "0000000010",  -- +0.0737
        4 => "1111100101",  -- -0.8591
        5 => "1111001011",  -- -1.6505
        6 => "1111111110",  -- -0.0676
        7 => "1111011110",  -- -1.0569
        8 => "1110111111",  -- -2.0179
        9 => "1111110001",  -- -0.4633
        10 => "1111010100",  -- -1.3678
        11 => "1111000111",  -- -1.7918
        12 => "0000000111",  -- +0.2150
        13 => "1111110110",  -- -0.3220
        14 => "1111111010",  -- -0.1807
        15 => "0000001110",  -- +0.4411
        16 => "0000001010",  -- +0.2998
        17 => "0000001111",  -- +0.4694
        18 => "0000010000",  -- +0.4977
        19 => "0000001010",  -- +0.3281
        20 => "0000001010",  -- +0.2998
        21 => "1111110101",  -- -0.3503
        22 => "1111101101",  -- -0.6047
        23 => "1111101000",  -- -0.7460
        24 => "1111101101",  -- -0.6047
        25 => "1111100000",  -- -1.0004
        26 => "1111011001",  -- -1.2265
        27 => "1111110111",  -- -0.2938
        28 => "1111100110",  -- -0.8025
        29 => "1111011100",  -- -1.1134
        30 => "0000000001",  -- +0.0454
        31 => "1111101110",  -- -0.5481
        32 => "1111100010",  -- -0.9439
        33 => "0000010011",  -- +0.5825
        34 => "0000000000",  -- -0.0111
        35 => "1111101110",  -- -0.5764
        36 => "0000011011",  -- +0.8368
        37 => "0000000111",  -- +0.2150
        38 => "1111110001",  -- -0.4633
        39 => "0000011010",  -- +0.8086
        40 => "0000000001",  -- +0.0454
        41 => "1111110000",  -- -0.4916
        42 => "0000001010",  -- +0.2998
        43 => "1111110010",  -- -0.4351
        44 => "1111100101",  -- -0.8591
        45 => "1111101000",  -- -0.7460
        46 => "1111010101",  -- -1.3396
        47 => "1111001010",  -- -1.6787
        48 => "1111010110",  -- -1.3113
        49 => "1111001011",  -- -1.6505
        50 => "1110111111",  -- -2.0179
        51 => "0000000100",  -- +0.1302
        52 => "0000000000",  -- -0.0111
        53 => "1111110010",  -- -0.4351
        54 => "0000100111",  -- +1.2326
        55 => "0000100011",  -- +1.0912
        56 => "0000001110",  -- +0.4411
        57 => "0000101111",  -- +1.4587
        58 => "0000100111",  -- +1.2043
        59 => "0000001100",  -- +0.3846
        60 => "0000110000",  -- +1.5152
        61 => "0000100110",  -- +1.1760
        62 => "0000001010",  -- +0.3281
        63 => "0000101101",  -- +1.4021
        64 => "0000011110",  -- +0.9499
        65 => "0000000110",  -- +0.1867
        66 => "0000101101",  -- +1.4021
        67 => "0000011001",  -- +0.7803
        68 => "0000000001",  -- +0.0172
        69 => "0000101101",  -- +1.4021
        70 => "0000010101",  -- +0.6673
        71 => "1111111101",  -- -0.0959
        72 => "1110010101",  -- -3.3464
        73 => "1110001011",  -- -3.6573
        74 => "1110001000",  -- -3.7421
        75 => "1111101010",  -- -0.6895
        76 => "1111010001",  -- -1.4809
        77 => "1110111001",  -- -2.2158
        78 => "1111111101",  -- -0.0959
        79 => "1111011110",  -- -1.0569
        80 => "1110111111",  -- -2.0462
        81 => "1111110100",  -- -0.3786
        82 => "1111010101",  -- -1.3396
        83 => "1111000101",  -- -1.8483
        84 => "0000000001",  -- +0.0454
        85 => "1111101101",  -- -0.6047
        86 => "1111110000",  -- -0.4916
        87 => "0000011000",  -- +0.7520
        88 => "0000010000",  -- +0.4977
        89 => "0000010111",  -- +0.7238
        90 => "0000011101",  -- +0.9216
        91 => "0000011001",  -- +0.7803
        92 => "0000011101",  -- +0.8934
        93 => "1111111111",  -- -0.0394
        94 => "1111111000",  -- -0.2655
        95 => "1111111000",  -- -0.2372
        96 => "1111011110",  -- -1.0569
        97 => "1111010011",  -- -1.3961
        98 => "1111010010",  -- -1.4526
        99 => "1111011010",  -- -1.1982
        100 => "1111001010",  -- -1.6787
        101 => "1111000101",  -- -1.8483
        102 => "1111011100",  -- -1.1134
        103 => "1111001001",  -- -1.7070
        104 => "1111000001",  -- -1.9614
        105 => "1111110001",  -- -0.4633
        106 => "1111100000",  -- -1.0004
        107 => "1111010011",  -- -1.3961
        108 => "1111111110",  -- -0.0676
        109 => "1111101101",  -- -0.6047
        110 => "1111011110",  -- -1.0569
        111 => "1111111110",  -- -0.0676
        112 => "1111101010",  -- -0.6895
        113 => "1111011111",  -- -1.0286
        114 => "1111101110",  -- -0.5481
        115 => "1111011101",  -- -1.0852
        116 => "1111010100",  -- -1.3678
        117 => "1111101010",  -- -0.6895
        118 => "1111100000",  -- -1.0004
        119 => "1111010111",  -- -1.2830
        120 => "1111101110",  -- -0.5764
        121 => "1111101010",  -- -0.6895
        122 => "1111100000",  -- -1.0004
        123 => "0000001101",  -- +0.4129
        124 => "0000001110",  -- +0.4411
        125 => "0000000000",  -- -0.0111
        126 => "0000010011",  -- +0.5825
        127 => "0000010100",  -- +0.6390
        128 => "1111111111",  -- -0.0394
        129 => "0000011110",  -- +0.9499
        130 => "0000011101",  -- +0.8934
        131 => "0000000010",  -- +0.0737
        132 => "0000101000",  -- +1.2608
        133 => "0000100100",  -- +1.1195
        134 => "0000001010",  -- +0.2998
        135 => "0000101101",  -- +1.4021
        136 => "0000100110",  -- +1.1760
        137 => "0000001110",  -- +0.4411
        138 => "0000101001",  -- +1.2891
        139 => "0000100001",  -- +1.0347
        140 => "0000001010",  -- +0.3281
        141 => "0000101111",  -- +1.4587
        142 => "0000100110",  -- +1.1760
        143 => "0000001110",  -- +0.4411
        144 => "1110001010",  -- -3.6856
        145 => "1110000100",  -- -3.8834
        146 => "1110000011",  -- -3.9117
        147 => "1111011010",  -- -1.1982
        148 => "1111001111",  -- -1.5374
        149 => "1110111100",  -- -2.1310
        150 => "0000001011",  -- +0.3563
        151 => "1111111010",  -- -0.1807
        152 => "1111011100",  -- -1.1134
        153 => "0000000011",  -- +0.1020
        154 => "1111101110",  -- -0.5481
        155 => "1111011000",  -- -1.2548
        156 => "0000000001",  -- +0.0454
        157 => "1111110001",  -- -0.4633
        158 => "1111101110",  -- -0.5764
        159 => "0000011011",  -- +0.8368
        160 => "0000010001",  -- +0.5259
        161 => "0000011001",  -- +0.7803
        162 => "0000011111",  -- +0.9782
        163 => "0000011000",  -- +0.7520
        164 => "0000011101",  -- +0.8934
        165 => "0000001010",  -- +0.3281
        166 => "0000000010",  -- +0.0737
        167 => "0000000011",  -- +0.1020
        168 => "1111100110",  -- -0.8025
        169 => "1111011100",  -- -1.1134
        170 => "1111011011",  -- -1.1700
        171 => "1111001111",  -- -1.5374
        172 => "1111000001",  -- -1.9614
        173 => "1110111110",  -- -2.0745
        174 => "1111010111",  -- -1.2830
        175 => "1111001000",  -- -1.7635
        176 => "1111000010",  -- -1.9331
        177 => "1111011110",  -- -1.0569
        178 => "1111001111",  -- -1.5374
        179 => "1111001000",  -- -1.7353
        180 => "1111010100",  -- -1.3678
        181 => "1111000111",  -- -1.7918
        182 => "1110111111",  -- -2.0179
        183 => "1111100001",  -- -0.9721
        184 => "1111010010",  -- -1.4526
        185 => "1111001011",  -- -1.6505
        186 => "1111010111",  -- -1.2830
        187 => "1111001001",  -- -1.7070
        188 => "1111000100",  -- -1.8766
        189 => "1111100111",  -- -0.7743
        190 => "1111011100",  -- -1.1134
        191 => "1111010111",  -- -1.2830
        192 => "0000010000",  -- +0.4977
        193 => "0000001010",  -- +0.2998
        194 => "0000000100",  -- +0.1302
        195 => "0000100000",  -- +1.0064
        196 => "0000011111",  -- +0.9782
        197 => "0000010110",  -- +0.6955
        198 => "0000010101",  -- +0.6673
        199 => "0000010110",  -- +0.6955
        200 => "0000000010",  -- +0.0737
        201 => "0000011110",  -- +0.9499
        202 => "0000011011",  -- +0.8368
        203 => "0000001000",  -- +0.2433
        204 => "0000101011",  -- +1.3456
        205 => "0000100011",  -- +1.0912
        206 => "0000011001",  -- +0.7803
        207 => "0000101110",  -- +1.4304
        208 => "0000100100",  -- +1.1195
        209 => "0000011010",  -- +0.8086
        210 => "0000101011",  -- +1.3456
        211 => "0000100110",  -- +1.1760
        212 => "0000011011",  -- +0.8368
        213 => "0000101111",  -- +1.4587
        214 => "0000101011",  -- +1.3456
        215 => "0000011111",  -- +0.9782
        216 => "1111000011",  -- -1.9049
        217 => "1110111111",  -- -2.0179
        218 => "1110111000",  -- -2.2440
        219 => "0000000111",  -- +0.2150
        220 => "0000000110",  -- +0.1867
        221 => "1111110100",  -- -0.3786
        222 => "0000010111",  -- +0.7238
        223 => "0000010001",  -- +0.5259
        224 => "1111110101",  -- -0.3503
        225 => "0000000001",  -- +0.0172
        226 => "1111110110",  -- -0.3220
        227 => "1111011011",  -- -1.1700
        228 => "1111111100",  -- -0.1242
        229 => "1111101111",  -- -0.5199
        230 => "1111100111",  -- -0.7743
        231 => "0000010110",  -- +0.6955
        232 => "0000001100",  -- +0.3846
        233 => "0000010100",  -- +0.6390
        234 => "0000011100",  -- +0.8651
        235 => "0000010100",  -- +0.6107
        236 => "0000010111",  -- +0.7238
        237 => "0000011001",  -- +0.7803
        238 => "0000010001",  -- +0.5259
        239 => "0000010000",  -- +0.4977
        240 => "0000000110",  -- +0.1867
        241 => "1111111101",  -- -0.0959
        242 => "1111111100",  -- -0.1242
        243 => "1111101100",  -- -0.6329
        244 => "1111100000",  -- -1.0004
        245 => "1111011101",  -- -1.0852
        246 => "1111101001",  -- -0.7177
        247 => "1111011101",  -- -1.0852
        248 => "1111011000",  -- -1.2548
        249 => "1111100000",  -- -1.0004
        250 => "1111010011",  -- -1.3961
        251 => "1111001111",  -- -1.5374
        252 => "1111001000",  -- -1.7353
        253 => "1110111100",  -- -2.1310
        254 => "1110111000",  -- -2.2440
        255 => "1111010110",  -- -1.3113
        256 => "1111001001",  -- -1.7070
        257 => "1111000110",  -- -1.8201
        258 => "1111010111",  -- -1.2830
        259 => "1111001010",  -- -1.6787
        260 => "1111000111",  -- -1.7918
        261 => "1111100110",  -- -0.8025
        262 => "1111011001",  -- -1.2265
        263 => "1111010110",  -- -1.3113
        264 => "0000010110",  -- +0.6955
        265 => "0000001011",  -- +0.3563
        266 => "0000001001",  -- +0.2715
        267 => "0000100110",  -- +1.1760
        268 => "0000100001",  -- +1.0347
        269 => "0000011100",  -- +0.8651
        270 => "0000010100",  -- +0.6107
        271 => "0000010010",  -- +0.5542
        272 => "1111111110",  -- -0.0676
        273 => "0000101001",  -- +1.2891
        274 => "0000100011",  -- +1.0912
        275 => "0000010100",  -- +0.6107
        276 => "0001000011",  -- +2.1088
        277 => "0000111001",  -- +1.7696
        278 => "0000110111",  -- +1.7131
        279 => "0000111111",  -- +1.9674
        280 => "0000110011",  -- +1.6000
        281 => "0000101111",  -- +1.4587
        282 => "0001000001",  -- +2.0240
        283 => "0000111010",  -- +1.7979
        284 => "0000110011",  -- +1.6000
        285 => "0000111010",  -- +1.8261
        286 => "0000110111",  -- +1.7131
        287 => "0000101110",  -- +1.4304
        288 => "0000001001",  -- +0.2715
        289 => "0000000111",  -- +0.2150
        290 => "1111110101",  -- -0.3503
        291 => "0000010100",  -- +0.6390
        292 => "0000010100",  -- +0.6107
        293 => "0000000000",  -- -0.0111
        294 => "0000010100",  -- +0.6390
        295 => "0000001110",  -- +0.4411
        296 => "1111110011",  -- -0.4068
        297 => "1111111001",  -- -0.2090
        298 => "1111101110",  -- -0.5764
        299 => "1111010100",  -- -1.3678
        300 => "1111100001",  -- -0.9721
        301 => "1111010101",  -- -1.3396
        302 => "1111001101",  -- -1.5939
        303 => "0000000101",  -- +0.1585
        304 => "1111111010",  -- -0.1807
        305 => "0000000001",  -- +0.0172
        306 => "0000011011",  -- +0.8368
        307 => "0000010011",  -- +0.5825
        308 => "0000010101",  -- +0.6673
        309 => "0000011101",  -- +0.9216
        310 => "0000010110",  -- +0.6955
        311 => "0000010101",  -- +0.6673
        312 => "0000011000",  -- +0.7520
        313 => "0000001111",  -- +0.4694
        314 => "0000001110",  -- +0.4411
        315 => "0000010000",  -- +0.4977
        316 => "0000000101",  -- +0.1585
        317 => "0000000010",  -- +0.0737
        318 => "0000000000",  -- -0.0111
        319 => "1111110100",  -- -0.3786
        320 => "1111101110",  -- -0.5481
        321 => "1111101101",  -- -0.6047
        322 => "1111011111",  -- -1.0286
        323 => "1111011011",  -- -1.1417
        324 => "1111011101",  -- -1.0852
        325 => "1111010001",  -- -1.4809
        326 => "1111001110",  -- -1.5657
        327 => "1111011101",  -- -1.0852
        328 => "1111010001",  -- -1.4809
        329 => "1111001110",  -- -1.5657
        330 => "1111100001",  -- -0.9721
        331 => "1111010100",  -- -1.3678
        332 => "1111010010",  -- -1.4526
        333 => "1111101000",  -- -0.7460
        334 => "1111011011",  -- -1.1417
        335 => "1111011001",  -- -1.2265
        336 => "0000001001",  -- +0.2715
        337 => "1111111111",  -- -0.0394
        338 => "1111111100",  -- -0.1242
        339 => "0000011110",  -- +0.9499
        340 => "0000011011",  -- +0.8368
        341 => "0000010010",  -- +0.5542
        342 => "0000010100",  -- +0.6107
        343 => "0000010011",  -- +0.5825
        344 => "1111111011",  -- -0.1524
        345 => "0000110000",  -- +1.4869
        346 => "0000101100",  -- +1.3739
        347 => "0000010111",  -- +0.7238
        348 => "0001000011",  -- +2.0805
        349 => "0000111011",  -- +1.8544
        350 => "0000110010",  -- +1.5717
        351 => "0000111101",  -- +1.9109
        352 => "0000110101",  -- +1.6565
        353 => "0000101001",  -- +1.2891
        354 => "0000111010",  -- +1.8261
        355 => "0000110110",  -- +1.6848
        356 => "0000100100",  -- +1.1195
        357 => "0000101001",  -- +1.2891
        358 => "0000100111",  -- +1.2326
        359 => "0000010010",  -- +0.5542
        360 => "0000010111",  -- +0.7238
        361 => "0000010101",  -- +0.6673
        362 => "0000000000",  -- -0.0111
        363 => "0000011001",  -- +0.7803
        364 => "0000011000",  -- +0.7520
        365 => "0000000001",  -- +0.0454
        366 => "0000011011",  -- +0.8368
        367 => "0000010100",  -- +0.6390
        368 => "1111111000",  -- -0.2372
        369 => "1111110111",  -- -0.2938
        370 => "1111101011",  -- -0.6612
        371 => "1111010010",  -- -1.4244
        372 => "1111011100",  -- -1.1134
        373 => "1111010001",  -- -1.4809
        374 => "1111000111",  -- -1.7918
        375 => "1111111100",  -- -0.1242
        376 => "1111110010",  -- -0.4351
        377 => "1111110101",  -- -0.3503
        378 => "0000010000",  -- +0.4977
        379 => "0000001001",  -- +0.2715
        380 => "0000001010",  -- +0.3281
        381 => "0000010101",  -- +0.6673
        382 => "0000001101",  -- +0.4129
        383 => "0000001100",  -- +0.3846
        384 => "0000010111",  -- +0.7238
        385 => "0000001110",  -- +0.4411
        386 => "0000001101",  -- +0.4129
        387 => "0000011001",  -- +0.7803
        388 => "0000001101",  -- +0.4129
        389 => "0000001011",  -- +0.3563
        390 => "0000001010",  -- +0.2998
        391 => "1111111101",  -- -0.0959
        392 => "1111111000",  -- -0.2372
        393 => "1111110001",  -- -0.4633
        394 => "1111100101",  -- -0.8308
        395 => "1111100011",  -- -0.9156
        396 => "1111010000",  -- -1.5092
        397 => "1111000101",  -- -1.8483
        398 => "1111000011",  -- -1.9049
        399 => "1111011101",  -- -1.0852
        400 => "1111010011",  -- -1.3961
        401 => "1111010010",  -- -1.4526
        402 => "1111011111",  -- -1.0286
        403 => "1111010100",  -- -1.3678
        404 => "1111010010",  -- -1.4244
        405 => "1111100010",  -- -0.9439
        406 => "1111011000",  -- -1.2548
        407 => "1111010110",  -- -1.3113
        408 => "0000000010",  -- +0.0737
        409 => "1111111001",  -- -0.2090
        410 => "1111111000",  -- -0.2655
        411 => "0000011000",  -- +0.7520
        412 => "0000010100",  -- +0.6107
        413 => "0000001010",  -- +0.2998
        414 => "0000100101",  -- +1.1478
        415 => "0000100101",  -- +1.1478
        416 => "0000001010",  -- +0.2998
        417 => "0000111100",  -- +1.8827
        418 => "0000111011",  -- +1.8544
        419 => "0000100001",  -- +1.0347
        420 => "0000111110",  -- +1.9392
        421 => "0000111010",  -- +1.8261
        422 => "0000101100",  -- +1.3739
        423 => "0001000010",  -- +2.0522
        424 => "0000111101",  -- +1.9109
        425 => "0000101010",  -- +1.3174
        426 => "0000111101",  -- +1.9109
        427 => "0000111100",  -- +1.8827
        428 => "0000100000",  -- +1.0064
        429 => "0000011110",  -- +0.9499
        430 => "0000100000",  -- +1.0064
        431 => "0000000000",  -- -0.0111
        432 => "0000011101",  -- +0.9216
        433 => "0000011100",  -- +0.8651
        434 => "0000000111",  -- +0.2150
        435 => "0000100010",  -- +1.0630
        436 => "0000100010",  -- +1.0630
        437 => "0000001000",  -- +0.2433
        438 => "0000011011",  -- +0.8368
        439 => "0000010101",  -- +0.6673
        440 => "1111111001",  -- -0.2090
        441 => "1111110001",  -- -0.4633
        442 => "1111100101",  -- -0.8308
        443 => "1111001110",  -- -1.5657
        444 => "1111101111",  -- -0.5199
        445 => "1111100100",  -- -0.8873
        446 => "1111011000",  -- -1.2548
        447 => "0000000111",  -- +0.2150
        448 => "1111111110",  -- -0.0676
        449 => "1111111101",  -- -0.0959
        450 => "0000001111",  -- +0.4694
        451 => "0000001000",  -- +0.2433
        452 => "0000001001",  -- +0.2715
        453 => "0000010100",  -- +0.6107
        454 => "0000001100",  -- +0.3846
        455 => "0000001011",  -- +0.3563
        456 => "0000010111",  -- +0.7238
        457 => "0000001111",  -- +0.4694
        458 => "0000001101",  -- +0.4129
        459 => "0000010010",  -- +0.5542
        460 => "0000000111",  -- +0.2150
        461 => "0000000100",  -- +0.1302
        462 => "0000000001",  -- +0.0172
        463 => "1111110100",  -- -0.3786
        464 => "1111101111",  -- -0.5199
        465 => "1111100100",  -- -0.8873
        466 => "1111011001",  -- -1.2265
        467 => "1111010110",  -- -1.3113
        468 => "1111010010",  -- -1.4244
        469 => "1111001001",  -- -1.7070
        470 => "1111001000",  -- -1.7353
        471 => "1111011100",  -- -1.1134
        472 => "1111010011",  -- -1.3961
        473 => "1111010010",  -- -1.4526
        474 => "1111011100",  -- -1.1134
        475 => "1111010100",  -- -1.3678
        476 => "1111010010",  -- -1.4244
        477 => "1111011101",  -- -1.0852
        478 => "1111010101",  -- -1.3396
        479 => "1111010011",  -- -1.3961
        480 => "0000000000",  -- -0.0111
        481 => "1111111000",  -- -0.2655
        482 => "1111110110",  -- -0.3220
        483 => "0000001100",  -- +0.3846
        484 => "0000001000",  -- +0.2433
        485 => "1111111111",  -- -0.0394
        486 => "0000100010",  -- +1.0630
        487 => "0000100010",  -- +1.0630
        488 => "0000000111",  -- +0.2150
        489 => "0001000010",  -- +2.0522
        490 => "0001000010",  -- +2.0522
        491 => "0000100110",  -- +1.1760
        492 => "0001000100",  -- +2.1370
        493 => "0001000100",  -- +2.1370
        494 => "0000110001",  -- +1.5435
        495 => "0001000100",  -- +2.1370
        496 => "0001000101",  -- +2.1653
        497 => "0000101100",  -- +1.3739
        498 => "0001000000",  -- +1.9957
        499 => "0001000011",  -- +2.1088
        500 => "0000100010",  -- +1.0630
        501 => "0000100011",  -- +1.0912
        502 => "0000101000",  -- +1.2608
        503 => "0000000001",  -- +0.0454
        504 => "0000100000",  -- +1.0064
        505 => "0000011110",  -- +0.9499
        506 => "0000001000",  -- +0.2433
        507 => "0000100101",  -- +1.1478
        508 => "0000100110",  -- +1.1760
        509 => "0000001000",  -- +0.2433
        510 => "0000011000",  -- +0.7520
        511 => "0000010011",  -- +0.5825
        512 => "1111110111",  -- -0.2938
        513 => "1111111001",  -- -0.2090
        514 => "1111101101",  -- -0.6047
        515 => "1111010111",  -- -1.2830
        516 => "0000000001",  -- +0.0172
        517 => "1111110101",  -- -0.3503
        518 => "1111101000",  -- -0.7460
        519 => "0000010101",  -- +0.6673
        520 => "0000001101",  -- +0.4129
        521 => "0000001001",  -- +0.2715
        522 => "0000010111",  -- +0.7238
        523 => "0000010000",  -- +0.4977
        524 => "0000010000",  -- +0.4977
        525 => "0000010101",  -- +0.6673
        526 => "0000001110",  -- +0.4411
        527 => "0000001101",  -- +0.4129
        528 => "0000010111",  -- +0.7238
        529 => "0000001110",  -- +0.4411
        530 => "0000001101",  -- +0.4129
        531 => "0000000100",  -- +0.1302
        532 => "1111111000",  -- -0.2372
        533 => "1111110111",  -- -0.2938
        534 => "1111101101",  -- -0.6047
        535 => "1111100000",  -- -1.0004
        536 => "1111011011",  -- -1.1417
        537 => "1111010100",  -- -1.3678
        538 => "1111001001",  -- -1.7070
        539 => "1111000111",  -- -1.7918
        540 => "1111011001",  -- -1.2265
        541 => "1111010001",  -- -1.4809
        542 => "1111010001",  -- -1.4809
        543 => "1111101001",  -- -0.7177
        544 => "1111100001",  -- -0.9721
        545 => "1111100000",  -- -1.0004
        546 => "1111100001",  -- -0.9721
        547 => "1111011001",  -- -1.2265
        548 => "1111011000",  -- -1.2548
        549 => "1111100011",  -- -0.9156
        550 => "1111011011",  -- -1.1700
        551 => "1111011010",  -- -1.1982
        552 => "0000000000",  -- -0.0111
        553 => "1111111000",  -- -0.2655
        554 => "1111111000",  -- -0.2372
        555 => "0000001000",  -- +0.2433
        556 => "0000000010",  -- +0.0737
        557 => "1111111101",  -- -0.0959
        558 => "0000010101",  -- +0.6673
        559 => "0000010100",  -- +0.6107
        560 => "1111111100",  -- -0.1242
        561 => "0000111100",  -- +1.8827
        562 => "0000111101",  -- +1.9109
        563 => "0000100011",  -- +1.0912
        564 => "0001000100",  -- +2.1370
        565 => "0001000111",  -- +2.2218
        566 => "0000110011",  -- +1.6000
        567 => "0001000011",  -- +2.0805
        568 => "0001000111",  -- +2.2218
        569 => "0000101101",  -- +1.4021
        570 => "0000111110",  -- +1.9392
        571 => "0001000011",  -- +2.1088
        572 => "0000100010",  -- +1.0630
        573 => "0000101011",  -- +1.3456
        574 => "0000110001",  -- +1.5435
        575 => "0000001100",  -- +0.3846
        576 => "0000011011",  -- +0.8368
        577 => "0000011010",  -- +0.8086
        578 => "1111111110",  -- -0.0676
        579 => "0000011101",  -- +0.8934
        580 => "0000011100",  -- +0.8651
        581 => "1111111101",  -- -0.0959
        582 => "0000010101",  -- +0.6673
        583 => "0000001110",  -- +0.4411
        584 => "1111110011",  -- -0.4068
        585 => "0000001011",  -- +0.3563
        586 => "1111111110",  -- -0.0676
        587 => "1111101010",  -- -0.6895
        588 => "0000000100",  -- +0.1302
        589 => "1111111000",  -- -0.2372
        590 => "1111101100",  -- -0.6329
        591 => "0000001010",  -- +0.3281
        592 => "0000000010",  -- +0.0737
        593 => "1111111100",  -- -0.1242
        594 => "0000001110",  -- +0.4411
        595 => "0000001000",  -- +0.2433
        596 => "0000000110",  -- +0.1867
        597 => "0000000101",  -- +0.1585
        598 => "1111111110",  -- -0.0676
        599 => "1111111101",  -- -0.0959
        600 => "0000000110",  -- +0.1867
        601 => "1111111101",  -- -0.0959
        602 => "1111111100",  -- -0.1242
        603 => "0000000110",  -- +0.1867
        604 => "1111111011",  -- -0.1524
        605 => "1111111000",  -- -0.2372
        606 => "1111110010",  -- -0.4351
        607 => "1111100101",  -- -0.8308
        608 => "1111100001",  -- -0.9721
        609 => "1111011111",  -- -1.0286
        610 => "1111010101",  -- -1.3396
        611 => "1111010011",  -- -1.3961
        612 => "1111101000",  -- -0.7460
        613 => "1111100001",  -- -0.9721
        614 => "1111100010",  -- -0.9439
        615 => "1111111111",  -- -0.0394
        616 => "1111111000",  -- -0.2372
        617 => "1111111000",  -- -0.2372
        618 => "1111101001",  -- -0.7177
        619 => "1111100011",  -- -0.9156
        620 => "1111100011",  -- -0.9156
        621 => "1111110100",  -- -0.3786
        622 => "1111101101",  -- -0.6047
        623 => "1111101101",  -- -0.6047
        624 => "0000000001",  -- +0.0454
        625 => "1111111010",  -- -0.1807
        626 => "1111111100",  -- -0.1242
        627 => "0000000100",  -- +0.1302
        628 => "1111111110",  -- -0.0676
        629 => "1111111100",  -- -0.1242
        630 => "0000010101",  -- +0.6673
        631 => "0000010100",  -- +0.6107
        632 => "0000000001",  -- +0.0172
        633 => "0000111001",  -- +1.7696
        634 => "0000111010",  -- +1.7979
        635 => "0000100010",  -- +1.0630
        636 => "0001000010",  -- +2.0522
        637 => "0001000101",  -- +2.1653
        638 => "0000110010",  -- +1.5717
        639 => "0001000011",  -- +2.0805
        640 => "0001001001",  -- +2.2784
        641 => "0000110000",  -- +1.4869
        642 => "0001000001",  -- +2.0240
        643 => "0001001000",  -- +2.2501
        644 => "0000101010",  -- +1.3174
        645 => "0000110111",  -- +1.7131
        646 => "0000111100",  -- +1.8827
        647 => "0000011101",  -- +0.8934
        648 => "0000011110",  -- +0.9499
        649 => "0000010111",  -- +0.7238
        650 => "1111111100",  -- -0.1242
        651 => "0000001011",  -- +0.3563
        652 => "0000000000",  -- -0.0111
        653 => "1111100100",  -- -0.8873
        654 => "0000001001",  -- +0.2715
        655 => "1111110110",  -- -0.3220
        656 => "1111011111",  -- -1.0286
        657 => "0000011111",  -- +0.9782
        658 => "0000010000",  -- +0.4977
        659 => "1111111101",  -- -0.0959
        660 => "0000000011",  -- +0.1020
        661 => "1111111010",  -- -0.1807
        662 => "1111101101",  -- -0.6047
        663 => "1111110100",  -- -0.3786
        664 => "1111101100",  -- -0.6329
        665 => "1111100100",  -- -0.8873
        666 => "1111101001",  -- -0.7177
        667 => "1111100011",  -- -0.9156
        668 => "1111100000",  -- -1.0004
        669 => "1111101001",  -- -0.7177
        670 => "1111100011",  -- -0.9156
        671 => "1111100001",  -- -0.9721
        672 => "0000000001",  -- +0.0172
        673 => "1111111010",  -- -0.1807
        674 => "1111111000",  -- -0.2372
        675 => "0000000001",  -- +0.0172
        676 => "1111111000",  -- -0.2655
        677 => "1111111000",  -- -0.2655
        678 => "1111101110",  -- -0.5764
        679 => "1111100101",  -- -0.8591
        680 => "1111100011",  -- -0.9156
        681 => "1111110110",  -- -0.3220
        682 => "1111101010",  -- -0.6895
        683 => "1111101101",  -- -0.6047
        684 => "0000000111",  -- +0.2150
        685 => "1111111101",  -- -0.0959
        686 => "0000000000",  -- -0.0111
        687 => "0000000001",  -- +0.0454
        688 => "1111111101",  -- -0.0959
        689 => "1111111011",  -- -0.1524
        690 => "1111110000",  -- -0.4916
        691 => "1111101111",  -- -0.5199
        692 => "1111101011",  -- -0.6612
        693 => "1111111101",  -- -0.0959
        694 => "1111111011",  -- -0.1524
        695 => "1111111000",  -- -0.2655
        696 => "1111111000",  -- -0.2655
        697 => "1111110011",  -- -0.4068
        698 => "1111110010",  -- -0.4351
        699 => "1111111001",  -- -0.2090
        700 => "1111110111",  -- -0.2938
        701 => "1111110010",  -- -0.4351
        702 => "0000011011",  -- +0.8368
        703 => "0000011001",  -- +0.7803
        704 => "0000001000",  -- +0.2433
        705 => "0000111001",  -- +1.7696
        706 => "0000110111",  -- +1.7131
        707 => "0000100000",  -- +1.0064
        708 => "0001000011",  -- +2.0805
        709 => "0001000011",  -- +2.1088
        710 => "0000101011",  -- +1.3456
        711 => "0001000011",  -- +2.0805
        712 => "0001001000",  -- +2.2501
        713 => "0000101100",  -- +1.3739
        714 => "0001000101",  -- +2.1653
        715 => "0001001010",  -- +2.3066
        716 => "0000110000",  -- +1.5152
        717 => "0001000011",  -- +2.1088
        718 => "0001000110",  -- +2.1936
        719 => "0000101110",  -- +1.4304
        720 => "0000100100",  -- +1.1195
        721 => "0000010101",  -- +0.6673
        722 => "0000000001",  -- +0.0172
        723 => "0000000010",  -- +0.0737
        724 => "1111101001",  -- -0.7177
        725 => "1111010101",  -- -1.3396
        726 => "1111111010",  -- -0.1807
        727 => "1111011010",  -- -1.1982
        728 => "1111001011",  -- -1.6505
        729 => "0000101011",  -- +1.3456
        730 => "0000010111",  -- +0.7238
        731 => "0000001010",  -- +0.2998
        732 => "0000010100",  -- +0.6107
        733 => "0000001100",  -- +0.3846
        734 => "1111111111",  -- -0.0394
        735 => "0000010001",  -- +0.5259
        736 => "0000001001",  -- +0.2715
        737 => "0000000000",  -- -0.0111
        738 => "0000000101",  -- +0.1585
        739 => "1111111111",  -- -0.0394
        740 => "1111111010",  -- -0.1807
        741 => "0000000100",  -- +0.1302
        742 => "0000000000",  -- -0.0111
        743 => "1111111100",  -- -0.1242
        744 => "0000010100",  -- +0.6390
        745 => "0000001111",  -- +0.4694
        746 => "0000001101",  -- +0.4129
        747 => "0000001001",  -- +0.2715
        748 => "0000000010",  -- +0.0737
        749 => "0000000011",  -- +0.1020
        750 => "1111100101",  -- -0.8591
        751 => "1111011110",  -- -1.0569
        752 => "1111100000",  -- -1.0004
        753 => "1111011011",  -- -1.1417
        754 => "1111010000",  -- -1.5092
        755 => "1111010101",  -- -1.3396
        756 => "0000001011",  -- +0.3563
        757 => "1111111110",  -- -0.0676
        758 => "0000000001",  -- +0.0454
        759 => "0000000110",  -- +0.1867
        760 => "0000000010",  -- +0.0737
        761 => "1111111100",  -- -0.1242
        762 => "1111110000",  -- -0.4916
        763 => "1111110010",  -- -0.4351
        764 => "1111100111",  -- -0.7743
        765 => "1111111001",  -- -0.2090
        766 => "1111111000",  -- -0.2655
        767 => "1111101111",  -- -0.5199
        768 => "0000000111",  -- +0.2150
        769 => "0000000011",  -- +0.1020
        770 => "1111111111",  -- -0.0394
        771 => "0000001000",  -- +0.2433
        772 => "0000000110",  -- +0.1867
        773 => "1111111101",  -- -0.0959
        774 => "0000010111",  -- +0.7238
        775 => "0000010100",  -- +0.6107
        776 => "0000000010",  -- +0.0737
        777 => "0000111110",  -- +1.9392
        778 => "0000111010",  -- +1.7979
        779 => "0000100001",  -- +1.0347
        780 => "0001000110",  -- +2.1936
        781 => "0001000011",  -- +2.1088
        782 => "0000100111",  -- +1.2326
        783 => "0001000011",  -- +2.1088
        784 => "0001000101",  -- +2.1653
        785 => "0000101001",  -- +1.2891
        786 => "0001000100",  -- +2.1370
        787 => "0001000110",  -- +2.1936
        788 => "0000101110",  -- +1.4304
        789 => "0001001100",  -- +2.3632
        790 => "0001001100",  -- +2.3632
        791 => "0000110111",  -- +1.7131
        792 => "0000100110",  -- +1.1760
        793 => "0000010100",  -- +0.6107
        794 => "0000000010",  -- +0.0737
        795 => "0000001100",  -- +0.3846
        796 => "1111101100",  -- -0.6329
        797 => "1111100000",  -- -1.0004
        798 => "1111110100",  -- -0.3786
        799 => "1111001110",  -- -1.5657
        800 => "1111000111",  -- -1.7918
        801 => "0000101101",  -- +1.4021
        802 => "0000010110",  -- +0.6955
        803 => "0000001110",  -- +0.4411
        804 => "0000100011",  -- +1.0912
        805 => "0000011101",  -- +0.8934
        806 => "0000010011",  -- +0.5825
        807 => "0000011011",  -- +0.8368
        808 => "0000010100",  -- +0.6390
        809 => "0000001101",  -- +0.4129
        810 => "0000011001",  -- +0.7803
        811 => "0000010100",  -- +0.6107
        812 => "0000001111",  -- +0.4694
        813 => "0000010000",  -- +0.4977
        814 => "0000001011",  -- +0.3563
        815 => "0000001000",  -- +0.2433
        816 => "0000000010",  -- +0.0737
        817 => "1111111101",  -- -0.0959
        818 => "1111111011",  -- -0.1524
        819 => "0000000101",  -- +0.1585
        820 => "0000000000",  -- -0.0111
        821 => "0000000001",  -- +0.0172
        822 => "1111111111",  -- -0.0394
        823 => "1111111001",  -- -0.2090
        824 => "1111111100",  -- -0.1242
        825 => "1111110010",  -- -0.4351
        826 => "1111100101",  -- -0.8591
        827 => "1111101000",  -- -0.7460
        828 => "1111111100",  -- -0.1242
        829 => "1111101101",  -- -0.6047
        830 => "1111101100",  -- -0.6329
        831 => "0000001111",  -- +0.4694
        832 => "0000001000",  -- +0.2433
        833 => "1111111110",  -- -0.0676
        834 => "1111111111",  -- -0.0394
        835 => "1111111011",  -- -0.1524
        836 => "1111101101",  -- -0.6047
        837 => "1111110010",  -- -0.4351
        838 => "1111101100",  -- -0.6329
        839 => "1111100001",  -- -0.9721
        840 => "0000010110",  -- +0.6955
        841 => "0000001111",  -- +0.4694
        842 => "0000000111",  -- +0.2150
        843 => "0000001100",  -- +0.3846
        844 => "0000001001",  -- +0.2715
        845 => "1111111110",  -- -0.0676
        846 => "0000000111",  -- +0.2150
        847 => "0000000001",  -- +0.0172
        848 => "1111110000",  -- -0.4916
        849 => "0000100001",  -- +1.0347
        850 => "0000011001",  -- +0.7803
        851 => "0000000001",  -- +0.0454
        852 => "0001000000",  -- +1.9957
        853 => "0000111010",  -- +1.8261
        854 => "0000011111",  -- +0.9782
        855 => "0001000100",  -- +2.1370
        856 => "0001000011",  -- +2.0805
        857 => "0000101000",  -- +1.2608
        858 => "0001000101",  -- +2.1653
        859 => "0001000110",  -- +2.1936
        860 => "0000101101",  -- +1.4021
        861 => "0001001000",  -- +2.2501
        862 => "0001001010",  -- +2.3066
        863 => "0000110000",  -- +1.5152
        864 => "0000011011",  -- +0.8368
        865 => "0000001000",  -- +0.2433
        866 => "1111111010",  -- -0.1807
        867 => "0000011010",  -- +0.8086
        868 => "1111110101",  -- -0.3503
        869 => "1111110001",  -- -0.4633
        870 => "1111110101",  -- -0.3503
        871 => "1111001100",  -- -1.6222
        872 => "1111001011",  -- -1.6505
        873 => "0000011100",  -- +0.8651
        874 => "0000000101",  -- +0.1585
        875 => "0000000001",  -- +0.0172
        876 => "0000101010",  -- +1.3174
        877 => "0000100101",  -- +1.1478
        878 => "0000011101",  -- +0.8934
        879 => "0000010110",  -- +0.6955
        880 => "0000010001",  -- +0.5259
        881 => "0000001100",  -- +0.3846
        882 => "0000000110",  -- +0.1867
        883 => "0000000001",  -- +0.0172
        884 => "1111111101",  -- -0.0959
        885 => "0000001110",  -- +0.4411
        886 => "0000001010",  -- +0.2998
        887 => "0000000110",  -- +0.1867
        888 => "0000000101",  -- +0.1585
        889 => "0000000001",  -- +0.0172
        890 => "1111111110",  -- -0.0676
        891 => "1111111010",  -- -0.1807
        892 => "1111110101",  -- -0.3503
        893 => "1111110110",  -- -0.3220
        894 => "0000000110",  -- +0.1867
        895 => "0000000000",  -- -0.0111
        896 => "0000000010",  -- +0.0737
        897 => "0000001010",  -- +0.2998
        898 => "1111111101",  -- -0.0959
        899 => "1111111111",  -- -0.0394
        900 => "1111011100",  -- -1.1134
        901 => "1111001100",  -- -1.6222
        902 => "1111001000",  -- -1.7635
        903 => "1111111101",  -- -0.0959
        904 => "1111110000",  -- -0.4916
        905 => "1111100100",  -- -0.8873
        906 => "0000010100",  -- +0.6107
        907 => "0000001001",  -- +0.2715
        908 => "1111111000",  -- -0.2372
        909 => "1111101110",  -- -0.5764
        910 => "1111100010",  -- -0.9439
        911 => "1111010100",  -- -1.3678
        912 => "0000000000",  -- -0.0111
        913 => "1111110100",  -- -0.3786
        914 => "1111101010",  -- -0.6895
        915 => "0000001011",  -- +0.3563
        916 => "0000000011",  -- +0.1020
        917 => "1111111000",  -- -0.2655
        918 => "1111110110",  -- -0.3220
        919 => "1111101011",  -- -0.6612
        920 => "1111011011",  -- -1.1700
        921 => "1111010011",  -- -1.3961
        922 => "1111000111",  -- -1.7918
        923 => "1110110001",  -- -2.4702
        924 => "1111110111",  -- -0.2938
        925 => "1111101100",  -- -0.6329
        926 => "1111010011",  -- -1.3961
        927 => "0000101011",  -- +1.3456
        928 => "0000100110",  -- +1.1760
        929 => "0000001110",  -- +0.4411
        930 => "0001000001",  -- +2.0240
        931 => "0001000000",  -- +1.9957
        932 => "0000100110",  -- +1.1760
        933 => "0000111101",  -- +1.9109
        934 => "0000111111",  -- +1.9674
        935 => "0000100010",  -- +1.0630
        936 => "0000001011",  -- +0.3563
        937 => "1111111100",  -- -0.1242
        938 => "1111101111",  -- -0.5199
        939 => "0000011111",  -- +0.9782
        940 => "0000000000",  -- -0.0111
        941 => "1111111110",  -- -0.0676
        942 => "0000010100",  -- +0.6390
        943 => "1111101111",  -- -0.5199
        944 => "1111110001",  -- -0.4633
        945 => "0000010000",  -- +0.4977
        946 => "1111111011",  -- -0.1524
        947 => "1111111000",  -- -0.2372
        948 => "0000100100",  -- +1.1195
        949 => "0000011111",  -- +0.9782
        950 => "0000011000",  -- +0.7520
        951 => "0000100111",  -- +1.2043
        952 => "0000100010",  -- +1.0630
        953 => "0000011101",  -- +0.8934
        954 => "0000100010",  -- +1.0630
        955 => "0000011101",  -- +0.9216
        956 => "0000011010",  -- +0.8086
        957 => "0000101010",  -- +1.3174
        958 => "0000100110",  -- +1.1760
        959 => "0000100010",  -- +1.0630
        960 => "0000010111",  -- +0.7238
        961 => "0000010011",  -- +0.5825
        962 => "0000010000",  -- +0.4977
        963 => "0000000110",  -- +0.1867
        964 => "0000000001",  -- +0.0172
        965 => "0000000001",  -- +0.0172
        966 => "0000001000",  -- +0.2433
        967 => "0000000010",  -- +0.0737
        968 => "0000000100",  -- +0.1302
        969 => "0000000101",  -- +0.1585
        970 => "1111111010",  -- -0.1807
        971 => "1111111011",  -- -0.1524
        972 => "1111011101",  -- -1.0852
        973 => "1111001110",  -- -1.5657
        974 => "1111000111",  -- -1.7918
        975 => "1111100101",  -- -0.8591
        976 => "1111010101",  -- -1.3396
        977 => "1111001000",  -- -1.7635
        978 => "0000010101",  -- +0.6673
        979 => "0000000101",  -- +0.1585
        980 => "1111110101",  -- -0.3503
        981 => "1111110011",  -- -0.4068
        982 => "1111100011",  -- -0.9156
        983 => "1111010100",  -- -1.3678
        984 => "1111111100",  -- -0.1242
        985 => "1111101110",  -- -0.5764
        986 => "1111100010",  -- -0.9439
        987 => "0000011101",  -- +0.9216
        988 => "0000010001",  -- +0.5259
        989 => "0000000101",  -- +0.1585
        990 => "0000000011",  -- +0.1020
        991 => "1111110101",  -- -0.3503
        992 => "1111100100",  -- -0.8873
        993 => "1111100011",  -- -0.9156
        994 => "1111010001",  -- -1.4809
        995 => "1110111100",  -- -2.1310
        996 => "1111010010",  -- -1.4526
        997 => "1111000001",  -- -1.9614
        998 => "1110101100",  -- -2.6115
        999 => "1111101011",  -- -0.6612
        1000 => "1111100000",  -- -1.0004
        1001 => "1111001101",  -- -1.5939
        1002 => "0000001111",  -- +0.4694
        1003 => "0000001010",  -- +0.2998
        1004 => "1111110010",  -- -0.4351
        1005 => "0000010111",  -- +0.7238
        1006 => "0000010011",  -- +0.5825
        1007 => "1111111000",  -- -0.2655
        1008 => "0000010000",  -- +0.4977
        1009 => "0000000111",  -- +0.2150
        1010 => "1111111000",  -- -0.2372
        1011 => "0000100000",  -- +1.0064
        1012 => "0000001100",  -- +0.3846
        1013 => "0000001000",  -- +0.2433
        1014 => "0000100111",  -- +1.2043
        1015 => "0000001010",  -- +0.3281
        1016 => "0000001001",  -- +0.2715
        1017 => "0000011000",  -- +0.7520
        1018 => "0000001001",  -- +0.2715
        1019 => "0000000010",  -- +0.0737
        1020 => "0000010101",  -- +0.6673
        1021 => "0000010100",  -- +0.6107
        1022 => "0000001001",  -- +0.2715
        1023 => "0000100111",  -- +1.2326
        1024 => "0000100100",  -- +1.1195
        1025 => "0000011011",  -- +0.8368
        1026 => "0000101110",  -- +1.4304
        1027 => "0000101000",  -- +1.2608
        1028 => "0000100100",  -- +1.1195
        1029 => "0000110101",  -- +1.6565
        1030 => "0000110000",  -- +1.5152
        1031 => "0000101101",  -- +1.4021
        1032 => "0000110100",  -- +1.6283
        1033 => "0000110000",  -- +1.4869
        1034 => "0000101101",  -- +1.4021
        1035 => "0000100000",  -- +1.0064
        1036 => "0000011011",  -- +0.8368
        1037 => "0000011100",  -- +0.8651
        1038 => "0000010100",  -- +0.6390
        1039 => "0000001111",  -- +0.4694
        1040 => "0000010010",  -- +0.5542
        1041 => "0000001010",  -- +0.3281
        1042 => "0000000011",  -- +0.1020
        1043 => "0000000010",  -- +0.0737
        1044 => "1111110001",  -- -0.4633
        1045 => "1111100110",  -- -0.8025
        1046 => "1111011111",  -- -1.0286
        1047 => "1111010110",  -- -1.3113
        1048 => "1111000110",  -- -1.8201
        1049 => "1110111010",  -- -2.1875
        1050 => "0000000001",  -- +0.0172
        1051 => "1111101111",  -- -0.5199
        1052 => "1111100001",  -- -0.9721
        1053 => "1111111000",  -- -0.2655
        1054 => "1111100111",  -- -0.7743
        1055 => "1111011011",  -- -1.1700
        1056 => "0000000000",  -- -0.0111
        1057 => "1111110001",  -- -0.4633
        1058 => "1111100110",  -- -0.8025
        1059 => "0000011000",  -- +0.7520
        1060 => "0000001001",  -- +0.2715
        1061 => "1111111011",  -- -0.1524
        1062 => "0000000010",  -- +0.0737
        1063 => "1111101110",  -- -0.5481
        1064 => "1111011110",  -- -1.0569
        1065 => "0000000100",  -- +0.1302
        1066 => "1111101110",  -- -0.5764
        1067 => "1111011011",  -- -1.1700
        1068 => "1111110100",  -- -0.3786
        1069 => "1111011111",  -- -1.0286
        1070 => "1111001101",  -- -1.5939
        1071 => "1111011111",  -- -1.0286
        1072 => "1111001110",  -- -1.5657
        1073 => "1110111111",  -- -2.0179
        1074 => "1111110011",  -- -0.4068
        1075 => "1111100101",  -- -0.8308
        1076 => "1111010011",  -- -1.3961
        1077 => "0000000001",  -- +0.0454
        1078 => "1111110110",  -- -0.3220
        1079 => "1111100000",  -- -1.0004
        1080 => "0000011011",  -- +0.8368
        1081 => "0000011000",  -- +0.7520
        1082 => "0000000111",  -- +0.2150
        1083 => "0000011111",  -- +0.9782
        1084 => "0000011000",  -- +0.7520
        1085 => "0000001110",  -- +0.4411
        1086 => "0000100110",  -- +1.1760
        1087 => "0000010100",  -- +0.6390
        1088 => "0000001101",  -- +0.4129
        1089 => "0000100111",  -- +1.2043
        1090 => "0000011101",  -- +0.9216
        1091 => "0000010011",  -- +0.5825
        1092 => "0000010001",  -- +0.5259
        1093 => "0000010001",  -- +0.5259
        1094 => "0000000010",  -- +0.0737
        1095 => "0000010100",  -- +0.6107
        1096 => "0000001111",  -- +0.4694
        1097 => "0000000010",  -- +0.0737
        1098 => "0000011011",  -- +0.8368
        1099 => "0000010101",  -- +0.6673
        1100 => "0000010000",  -- +0.4977
        1101 => "0000100001",  -- +1.0347
        1102 => "0000011101",  -- +0.8934
        1103 => "0000011000",  -- +0.7520
        1104 => "0000100110",  -- +1.1760
        1105 => "0000100000",  -- +1.0064
        1106 => "0000011110",  -- +0.9499
        1107 => "0000101001",  -- +1.2891
        1108 => "0000100101",  -- +1.1478
        1109 => "0000100101",  -- +1.1478
        1110 => "0000100100",  -- +1.1195
        1111 => "0000011101",  -- +0.9216
        1112 => "0000011111",  -- +0.9782
        1113 => "0000001100",  -- +0.3846
        1114 => "0000001001",  -- +0.2715
        1115 => "0000000111",  -- +0.2150
        1116 => "0000001010",  -- +0.2998
        1117 => "0000000011",  -- +0.1020
        1118 => "1111111101",  -- -0.0959
        1119 => "1111101111",  -- -0.5199
        1120 => "1111100011",  -- -0.9156
        1121 => "1111011000",  -- -1.2548
        1122 => "1111101101",  -- -0.6047
        1123 => "1111011011",  -- -1.1417
        1124 => "1111001111",  -- -1.5374
        1125 => "0000000111",  -- +0.2150
        1126 => "1111111000",  -- -0.2655
        1127 => "1111101100",  -- -0.6329
        1128 => "0000001110",  -- +0.4411
        1129 => "0000000001",  -- +0.0172
        1130 => "1111110111",  -- -0.2938
        1131 => "0000000110",  -- +0.1867
        1132 => "1111110101",  -- -0.3503
        1133 => "1111100111",  -- -0.7743
        1134 => "1111110110",  -- -0.3220
        1135 => "1111011111",  -- -1.0286
        1136 => "1111001111",  -- -1.5374
        1137 => "0000000011",  -- +0.1020
        1138 => "1111101010",  -- -0.6895
        1139 => "1111011000",  -- -1.2548
        1140 => "1111111100",  -- -0.1242
        1141 => "1111100101",  -- -0.8591
        1142 => "1111010100",  -- -1.3678
        1143 => "1111101110",  -- -0.5481
        1144 => "1111011011",  -- -1.1700
        1145 => "1111001110",  -- -1.5657
        1146 => "0000000001",  -- +0.0454
        1147 => "1111101110",  -- -0.5481
        1148 => "1111100010",  -- -0.9439
        1149 => "0000001011",  -- +0.3563
        1150 => "1111111000",  -- -0.2372
        1151 => "1111101001",  -- -0.7177
        1152 => "0000010101",  -- +0.6673
        1153 => "0000010101",  -- +0.6673
        1154 => "0000000011",  -- +0.1020
        1155 => "0000100000",  -- +1.0064
        1156 => "0000011101",  -- +0.8934
        1157 => "0000010001",  -- +0.5259
        1158 => "0000011110",  -- +0.9499
        1159 => "0000010100",  -- +0.6390
        1160 => "0000001001",  -- +0.2715
        1161 => "0000011111",  -- +0.9782
        1162 => "0000011000",  -- +0.7520
        1163 => "0000001010",  -- +0.2998
        1164 => "0000011111",  -- +0.9782
        1165 => "0000011100",  -- +0.8651
        1166 => "0000001011",  -- +0.3563
        1167 => "0000011001",  -- +0.7803
        1168 => "0000010011",  -- +0.5825
        1169 => "0000000100",  -- +0.1302
        1170 => "0000010111",  -- +0.7238
        1171 => "0000010100",  -- +0.6390
        1172 => "0000001010",  -- +0.2998
        1173 => "0000010110",  -- +0.6955
        1174 => "0000010001",  -- +0.5259
        1175 => "0000001001",  -- +0.2715
        1176 => "0000001010",  -- +0.2998
        1177 => "0000000011",  -- +0.1020
        1178 => "1111111101",  -- -0.0959
        1179 => "0000011100",  -- +0.8651
        1180 => "0000010111",  -- +0.7238
        1181 => "0000010011",  -- +0.5825
        1182 => "0000100100",  -- +1.1195
        1183 => "0000011100",  -- +0.8651
        1184 => "0000011001",  -- +0.7803
        1185 => "0000011101",  -- +0.8934
        1186 => "0000010101",  -- +0.6673
        1187 => "0000010100",  -- +0.6107
        1188 => "0000100111",  -- +1.2326
        1189 => "0000100100",  -- +1.1195
        1190 => "0000011110",  -- +0.9499
        1191 => "0000100000",  -- +1.0064
        1192 => "0000010101",  -- +0.6673
        1193 => "0000001101",  -- +0.4129
        1194 => "1111111111",  -- -0.0394
        1195 => "1111101110",  -- -0.5481
        1196 => "1111100100",  -- -0.8873
        1197 => "0000010010",  -- +0.5542
        1198 => "0000000001",  -- +0.0454
        1199 => "1111110111",  -- -0.2938
        1200 => "0000001001",  -- +0.2715
        1201 => "1111111001",  -- -0.2090
        1202 => "1111101110",  -- -0.5764
        1203 => "1111110101",  -- -0.3503
        1204 => "1111100011",  -- -0.9156
        1205 => "1111010101",  -- -1.3396
        1206 => "1111101110",  -- -0.5764
        1207 => "1111011000",  -- -1.2548
        1208 => "1111001000",  -- -1.7353
        1209 => "1111111111",  -- -0.0394
        1210 => "1111101000",  -- -0.7460
        1211 => "1111011001",  -- -1.2265
        1212 => "0000000000",  -- -0.0111
        1213 => "1111101001",  -- -0.7177
        1214 => "1111011100",  -- -1.1134
        1215 => "0000000011",  -- +0.1020
        1216 => "1111101111",  -- -0.5199
        1217 => "1111100101",  -- -0.8308
        1218 => "0000001101",  -- +0.4129
        1219 => "1111111000",  -- -0.2372
        1220 => "1111101110",  -- -0.5481
        1221 => "0000000111",  -- +0.2150
        1222 => "1111110010",  -- -0.4351
        1223 => "1111100101",  -- -0.8308
        1224 => "0000001010",  -- +0.3281
        1225 => "0000001010",  -- +0.3281
        1226 => "1111111000",  -- -0.2655
        1227 => "0000011101",  -- +0.9216
        1228 => "0000011001",  -- +0.7803
        1229 => "0000001110",  -- +0.4411
        1230 => "0000100101",  -- +1.1478
        1231 => "0000011101",  -- +0.9216
        1232 => "0000010010",  -- +0.5542
        1233 => "0000011101",  -- +0.9216
        1234 => "0000010100",  -- +0.6390
        1235 => "0000001000",  -- +0.2433
        1236 => "0000100110",  -- +1.1760
        1237 => "0000011100",  -- +0.8651
        1238 => "0000001111",  -- +0.4694
        1239 => "0000101011",  -- +1.3456
        1240 => "0000100010",  -- +1.0630
        1241 => "0000010101",  -- +0.6673
        1242 => "0000100111",  -- +1.2043
        1243 => "0000100110",  -- +1.1760
        1244 => "0000010110",  -- +0.6955
        1245 => "0000010001",  -- +0.5259
        1246 => "0000001010",  -- +0.2998
        1247 => "1111111101",  -- -0.0959
        1248 => "1111111010",  -- -0.1807
        1249 => "1111110001",  -- -0.4633
        1250 => "1111100110",  -- -0.8025
        1251 => "0000001101",  -- +0.4129
        1252 => "0000001010",  -- +0.3281
        1253 => "1111111111",  -- -0.0394
        1254 => "0000011010",  -- +0.8086
        1255 => "0000001101",  -- +0.4129
        1256 => "0000000101",  -- +0.1585
        1257 => "0000011000",  -- +0.7520
        1258 => "0000001100",  -- +0.3846
        1259 => "0000001001",  -- +0.2715
        1260 => "0000100000",  -- +1.0064
        1261 => "0000011011",  -- +0.8368
        1262 => "0000010110",  -- +0.6955
        1263 => "0000100100",  -- +1.1195
        1264 => "0000011010",  -- +0.8086
        1265 => "0000010011",  -- +0.5825
        1266 => "0000010100",  -- +0.6390
        1267 => "0000000110",  -- +0.1867
        1268 => "1111111011",  -- -0.1524
        1269 => "0000010000",  -- +0.4977
        1270 => "1111111110",  -- -0.0676
        1271 => "1111110000",  -- -0.4916
        1272 => "1111110101",  -- -0.3503
        1273 => "1111100010",  -- -0.9439
        1274 => "1111010011",  -- -1.3961
        1275 => "1111101001",  -- -0.7177
        1276 => "1111011001",  -- -1.2265
        1277 => "1111001001",  -- -1.7070
        1278 => "1111110101",  -- -0.3503
        1279 => "1111100101",  -- -0.8591
        1280 => "1111010110",  -- -1.3113
        1281 => "1111111111",  -- -0.0394
        1282 => "1111101110",  -- -0.5764
        1283 => "1111100001",  -- -0.9721
        1284 => "0000000100",  -- +0.1302
        1285 => "1111110011",  -- -0.4068
        1286 => "1111101001",  -- -0.7177
        1287 => "0000001010",  -- +0.3281
        1288 => "1111111010",  -- -0.1807
        1289 => "1111110000",  -- -0.4916
        1290 => "0000000101",  -- +0.1585
        1291 => "1111110011",  -- -0.4068
        1292 => "1111101000",  -- -0.7460
        1293 => "1111111000",  -- -0.2372
        1294 => "1111100110",  -- -0.8025
        1295 => "1111011010",  -- -1.1982
        1296 => "0000000001",  -- +0.0454
        1297 => "0000000010",  -- +0.0737
        1298 => "1111101110",  -- -0.5481
        1299 => "0000011011",  -- +0.8368
        1300 => "0000010101",  -- +0.6673
        1301 => "0000001011",  -- +0.3563
        1302 => "0000101110",  -- +1.4304
        1303 => "0000100111",  -- +1.2043
        1304 => "0000011101",  -- +0.8934
        1305 => "0000101101",  -- +1.4021
        1306 => "0000100100",  -- +1.1195
        1307 => "0000011011",  -- +0.8368
        1308 => "0000101011",  -- +1.3456
        1309 => "0000100000",  -- +1.0064
        1310 => "0000010111",  -- +0.7238
        1311 => "0000101101",  -- +1.4021
        1312 => "0000100011",  -- +1.0912
        1313 => "0000011001",  -- +0.7803
        1314 => "0000101000",  -- +1.2608
        1315 => "0000100100",  -- +1.1195
        1316 => "0000010110",  -- +0.6955
        1317 => "0000011001",  -- +0.7803
        1318 => "0000001011",  -- +0.3563
        1319 => "0000000001",  -- +0.0172
        1320 => "0000000010",  -- +0.0737
        1321 => "1111110110",  -- -0.3220
        1322 => "1111101100",  -- -0.6329
        1323 => "0000001010",  -- +0.3281
        1324 => "0000000110",  -- +0.1867
        1325 => "1111111000",  -- -0.2372
        1326 => "0000011001",  -- +0.7803
        1327 => "0000001011",  -- +0.3563
        1328 => "0000000001",  -- +0.0454
        1329 => "0000010101",  -- +0.6673
        1330 => "0000001000",  -- +0.2433
        1331 => "0000000010",  -- +0.0737
        1332 => "0000010100",  -- +0.6390
        1333 => "0000001101",  -- +0.4129
        1334 => "0000000111",  -- +0.2150
        1335 => "0000010110",  -- +0.6955
        1336 => "0000001100",  -- +0.3846
        1337 => "0000000100",  -- +0.1302
        1338 => "0000010110",  -- +0.6955
        1339 => "0000001000",  -- +0.2433
        1340 => "1111111100",  -- -0.1242
        1341 => "0000000010",  -- +0.0737
        1342 => "1111110000",  -- -0.4916
        1343 => "1111100010",  -- -0.9439
        1344 => "1111100000",  -- -1.0004
        1345 => "1111001101",  -- -1.5939
        1346 => "1110111101",  -- -2.1027
        1347 => "1111101001",  -- -0.7177
        1348 => "1111011010",  -- -1.1982
        1349 => "1111001010",  -- -1.6787
        1350 => "0000000000",  -- -0.0111
        1351 => "1111110000",  -- -0.4916
        1352 => "1111100010",  -- -0.9439
        1353 => "0000000010",  -- +0.0737
        1354 => "1111110010",  -- -0.4351
        1355 => "1111100110",  -- -0.8025
        1356 => "0000000010",  -- +0.0737
        1357 => "1111110010",  -- -0.4351
        1358 => "1111101000",  -- -0.7460
        1359 => "0000001010",  -- +0.3281
        1360 => "1111111010",  -- -0.1807
        1361 => "1111110001",  -- -0.4633
        1362 => "0000000101",  -- +0.1585
        1363 => "1111110100",  -- -0.3786
        1364 => "1111101001",  -- -0.7177
        1365 => "1111110111",  -- -0.2938
        1366 => "1111100101",  -- -0.8308
        1367 => "1111011001",  -- -1.2265
        1368 => "0000000001",  -- +0.0172
        1369 => "0000000010",  -- +0.0737
        1370 => "1111101010",  -- -0.6895
        1371 => "0000010111",  -- +0.7238
        1372 => "0000010011",  -- +0.5825
        1373 => "0000001000",  -- +0.2433
        1374 => "0000101100",  -- +1.3739
        1375 => "0000100111",  -- +1.2043
        1376 => "0000011110",  -- +0.9499
        1377 => "0000110001",  -- +1.5435
        1378 => "0000101001",  -- +1.2891
        1379 => "0000100100",  -- +1.1195
        1380 => "0000110010",  -- +1.5717
        1381 => "0000101000",  -- +1.2608
        1382 => "0000100011",  -- +1.0912
        1383 => "0000110001",  -- +1.5435
        1384 => "0000100111",  -- +1.2326
        1385 => "0000100000",  -- +1.0064
        1386 => "0000100111",  -- +1.2326
        1387 => "0000011101",  -- +0.8934
        1388 => "0000010100",  -- +0.6107
        1389 => "0000100010",  -- +1.0630
        1390 => "0000001101",  -- +0.4129
        1391 => "0000000111",  -- +0.2150
        1392 => "0000011000",  -- +0.7520
        1393 => "0000000110",  -- +0.1867
        1394 => "1111111110",  -- -0.0676
        1395 => "0000011000",  -- +0.7520
        1396 => "0000010001",  -- +0.5259
        1397 => "0000000011",  -- +0.1020
        1398 => "0000011110",  -- +0.9499
        1399 => "0000010001",  -- +0.5259
        1400 => "0000000110",  -- +0.1867
        1401 => "0000011100",  -- +0.8651
        1402 => "0000001100",  -- +0.3846
        1403 => "0000000100",  -- +0.1302
        1404 => "0000011100",  -- +0.8651
        1405 => "0000010001",  -- +0.5259
        1406 => "0000001010",  -- +0.2998
        1407 => "0000011010",  -- +0.8086
        1408 => "0000001101",  -- +0.4129
        1409 => "0000000011",  -- +0.1020
        1410 => "0000010011",  -- +0.5825
        1411 => "0000000011",  -- +0.1020
        1412 => "1111111000",  -- -0.2655
        1413 => "1111110011",  -- -0.4068
        1414 => "1111100001",  -- -0.9721
        1415 => "1111010010",  -- -1.4244
        1416 => "1111100010",  -- -0.9439
        1417 => "1111010000",  -- -1.5092
        1418 => "1111000000",  -- -1.9897
        1419 => "1111110101",  -- -0.3503
        1420 => "1111100101",  -- -0.8591
        1421 => "1111010101",  -- -1.3396
        1422 => "0000000011",  -- +0.1020
        1423 => "1111110100",  -- -0.3786
        1424 => "1111100101",  -- -0.8308
        1425 => "0000000000",  -- -0.0111
        1426 => "1111101111",  -- -0.5199
        1427 => "1111100100",  -- -0.8873
        1428 => "1111111111",  -- -0.0394
        1429 => "1111101110",  -- -0.5481
        1430 => "1111100101",  -- -0.8308
        1431 => "0000010100",  -- +0.6107
        1432 => "0000000011",  -- +0.1020
        1433 => "1111111010",  -- -0.1807
        1434 => "0000001010",  -- +0.2998
        1435 => "1111111000",  -- -0.2372
        1436 => "1111101101",  -- -0.6047
        1437 => "1111111110",  -- -0.0676
        1438 => "1111101101",  -- -0.6047
        1439 => "1111100000",  -- -1.0004
        1440 => "0000000111",  -- +0.2150
        1441 => "0000001010",  -- +0.3281
        1442 => "1111101101",  -- -0.6047
        1443 => "0000010101",  -- +0.6673
        1444 => "0000010100",  -- +0.6107
        1445 => "0000000010",  -- +0.0737
        1446 => "0000100111",  -- +1.2326
        1447 => "0000100100",  -- +1.1195
        1448 => "0000011100",  -- +0.8651
        1449 => "0000101001",  -- +1.2891
        1450 => "0000100010",  -- +1.0630
        1451 => "0000011111",  -- +0.9782
        1452 => "0000101010",  -- +1.3174
        1453 => "0000100010",  -- +1.0630
        1454 => "0000011101",  -- +0.9216
        1455 => "0000101100",  -- +1.3739
        1456 => "0000100010",  -- +1.0630
        1457 => "0000011011",  -- +0.8368
        1458 => "0000011100",  -- +0.8651
        1459 => "0000001001",  -- +0.2715
        1460 => "0000000011",  -- +0.1020
        1461 => "0000000011",  -- +0.1020
        1462 => "1111100101",  -- -0.8308
        1463 => "1111100100",  -- -0.8873
        1464 => "0000011000",  -- +0.7520
        1465 => "0000000000",  -- -0.0111
        1466 => "1111111010",  -- -0.1807
        1467 => "0000100011",  -- +1.0912
        1468 => "0000011001",  -- +0.7803
        1469 => "0000001011",  -- +0.3563
        1470 => "0000011110",  -- +0.9499
        1471 => "0000010010",  -- +0.5542
        1472 => "0000000011",  -- +0.1020
        1473 => "0000011110",  -- +0.9499
        1474 => "0000001101",  -- +0.4129
        1475 => "0000000010",  -- +0.0737
        1476 => "0000011101",  -- +0.9216
        1477 => "0000010000",  -- +0.4977
        1478 => "0000000101",  -- +0.1585
        1479 => "0000011011",  -- +0.8368
        1480 => "0000001100",  -- +0.3846
        1481 => "0000000001",  -- +0.0172
        1482 => "0000001001",  -- +0.2715
        1483 => "1111111000",  -- -0.2655
        1484 => "1111101011",  -- -0.6612
        1485 => "1111110000",  -- -0.4916
        1486 => "1111011110",  -- -1.0569
        1487 => "1111010001",  -- -1.4809
        1488 => "1111101011",  -- -0.6612
        1489 => "1111011010",  -- -1.1982
        1490 => "1111001010",  -- -1.6787
        1491 => "1111111000",  -- -0.2655
        1492 => "1111101000",  -- -0.7460
        1493 => "1111011001",  -- -1.2265
        1494 => "0000000000",  -- -0.0111
        1495 => "1111110000",  -- -0.4916
        1496 => "1111100010",  -- -0.9439
        1497 => "1111110111",  -- -0.2938
        1498 => "1111100111",  -- -0.7743
        1499 => "1111011011",  -- -1.1700
        1500 => "1111111000",  -- -0.2372
        1501 => "1111101000",  -- -0.7460
        1502 => "1111011110",  -- -1.0569
        1503 => "0000001100",  -- +0.3846
        1504 => "1111111100",  -- -0.1242
        1505 => "1111110011",  -- -0.4068
        1506 => "0000001000",  -- +0.2433
        1507 => "1111110111",  -- -0.2938
        1508 => "1111101100",  -- -0.6329
        1509 => "0000000001",  -- +0.0172
        1510 => "1111101111",  -- -0.5199
        1511 => "1111100011",  -- -0.9156
        1512 => "0000001100",  -- +0.3846
        1513 => "0000010010",  -- +0.5542
        1514 => "1111101110",  -- -0.5764
        1515 => "0000010011",  -- +0.5825
        1516 => "0000010100",  -- +0.6390
        1517 => "1111111011",  -- -0.1524
        1518 => "0000100101",  -- +1.1478
        1519 => "0000100011",  -- +1.0912
        1520 => "0000010110",  -- +0.6955
        1521 => "0000100111",  -- +1.2043
        1522 => "0000100001",  -- +1.0347
        1523 => "0000011101",  -- +0.9216
        1524 => "0000100010",  -- +1.0630
        1525 => "0000011100",  -- +0.8651
        1526 => "0000010101",  -- +0.6673
        1527 => "0000100011",  -- +1.0912
        1528 => "0000011010",  -- +0.8086
        1529 => "0000010000",  -- +0.4977
        1530 => "1111111001",  -- -0.2090
        1531 => "1111011111",  -- -1.0286
        1532 => "1111011101",  -- -1.0852
        1533 => "1111010111",  -- -1.2830
        1534 => "1110110001",  -- -2.4702
        1535 => "1110110011",  -- -2.4136
        1536 => "0000001001",  -- +0.2715
        1537 => "1111101100",  -- -0.6329
        1538 => "1111101000",  -- -0.7460
        1539 => "0000100101",  -- +1.1478
        1540 => "0000011000",  -- +0.7520
        1541 => "0000001010",  -- +0.3281
        1542 => "0000011100",  -- +0.8651
        1543 => "0000001111",  -- +0.4694
        1544 => "1111111111",  -- -0.0394
        1545 => "0000011000",  -- +0.7520
        1546 => "0000000110",  -- +0.1867
        1547 => "1111111000",  -- -0.2372
        1548 => "0000010111",  -- +0.7238
        1549 => "0000000110",  -- +0.1867
        1550 => "1111111000",  -- -0.2372
        1551 => "0000001111",  -- +0.4694
        1552 => "1111111110",  -- -0.0676
        1553 => "1111110000",  -- -0.4916
        1554 => "1111111111",  -- -0.0394
        1555 => "1111101110",  -- -0.5764
        1556 => "1111100000",  -- -1.0004
        1557 => "1111110000",  -- -0.4916
        1558 => "1111011111",  -- -1.0286
        1559 => "1111010010",  -- -1.4526
        1560 => "1111100110",  -- -0.8025
        1561 => "1111010101",  -- -1.3396
        1562 => "1111001000",  -- -1.7635
        1563 => "1111110110",  -- -0.3220
        1564 => "1111100110",  -- -0.8025
        1565 => "1111010111",  -- -1.2830
        1566 => "1111111001",  -- -0.2090
        1567 => "1111101010",  -- -0.6895
        1568 => "1111011011",  -- -1.1417
        1569 => "1111110011",  -- -0.4068
        1570 => "1111100100",  -- -0.8873
        1571 => "1111010111",  -- -1.2830
        1572 => "1111110101",  -- -0.3503
        1573 => "1111100101",  -- -0.8591
        1574 => "1111011011",  -- -1.1417
        1575 => "1111111001",  -- -0.2090
        1576 => "1111101001",  -- -0.7177
        1577 => "1111100000",  -- -1.0004
        1578 => "1111111000",  -- -0.2372
        1579 => "1111100111",  -- -0.7743
        1580 => "1111011100",  -- -1.1134
        1581 => "1111110101",  -- -0.3503
        1582 => "1111100100",  -- -0.8873
        1583 => "1111010111",  -- -1.2830
        1584 => "0000000110",  -- +0.1867
        1585 => "0000001100",  -- +0.3846
        1586 => "1111100010",  -- -0.9439
        1587 => "0000001010",  -- +0.2998
        1588 => "0000001110",  -- +0.4411
        1589 => "1111101101",  -- -0.6047
        1590 => "0000100010",  -- +1.0630
        1591 => "0000100010",  -- +1.0630
        1592 => "0000010001",  -- +0.5259
        1593 => "0000101010",  -- +1.3174
        1594 => "0000100110",  -- +1.1760
        1595 => "0000011111",  -- +0.9782
        1596 => "0000100110",  -- +1.1760
        1597 => "0000100001",  -- +1.0347
        1598 => "0000010110",  -- +0.6955
        1599 => "0000100000",  -- +1.0064
        1600 => "0000011000",  -- +0.7520
        1601 => "0000001010",  -- +0.2998
        1602 => "1111111101",  -- -0.0959
        1603 => "1111011101",  -- -1.0852
        1604 => "1111011110",  -- -1.0569
        1605 => "1111011111",  -- -1.0286
        1606 => "1110110010",  -- -2.4419
        1607 => "1110111000",  -- -2.2440
        1608 => "0000001011",  -- +0.3563
        1609 => "1111101001",  -- -0.7177
        1610 => "1111100111",  -- -0.7743
        1611 => "0000011111",  -- +0.9782
        1612 => "0000010001",  -- +0.5259
        1613 => "0000000100",  -- +0.1302
        1614 => "0000010010",  -- +0.5542
        1615 => "0000000011",  -- +0.1020
        1616 => "1111110010",  -- -0.4351
        1617 => "0000001101",  -- +0.4129
        1618 => "1111111010",  -- -0.1807
        1619 => "1111101011",  -- -0.6612
        1620 => "0000001101",  -- +0.4129
        1621 => "1111111010",  -- -0.1807
        1622 => "1111101100",  -- -0.6329
        1623 => "0000000001",  -- +0.0454
        1624 => "1111101111",  -- -0.5199
        1625 => "1111100000",  -- -1.0004
        1626 => "1111110111",  -- -0.2938
        1627 => "1111100101",  -- -0.8591
        1628 => "1111010111",  -- -1.2830
        1629 => "1111100110",  -- -0.8025
        1630 => "1111010101",  -- -1.3396
        1631 => "1111001000",  -- -1.7635
        1632 => "1111100010",  -- -0.9439
        1633 => "1111010001",  -- -1.4809
        1634 => "1111000011",  -- -1.9049
        1635 => "1111110011",  -- -0.4068
        1636 => "1111100011",  -- -0.9156
        1637 => "1111010100",  -- -1.3678
        1638 => "1111110100",  -- -0.3786
        1639 => "1111100101",  -- -0.8591
        1640 => "1111010110",  -- -1.3113
        1641 => "1111101011",  -- -0.6612
        1642 => "1111011011",  -- -1.1700
        1643 => "1111001110",  -- -1.5657
        1644 => "1111110001",  -- -0.4633
        1645 => "1111100001",  -- -0.9721
        1646 => "1111010111",  -- -1.2830
        1647 => "1111101000",  -- -0.7460
        1648 => "1111011000",  -- -1.2548
        1649 => "1111001111",  -- -1.5374
        1650 => "1111011111",  -- -1.0286
        1651 => "1111001110",  -- -1.5657
        1652 => "1111000011",  -- -1.9049
        1653 => "1111101000",  -- -0.7460
        1654 => "1111010111",  -- -1.2830
        1655 => "1111001010",  -- -1.6787
        1656 => "0000000001",  -- +0.0172
        1657 => "0000001000",  -- +0.2433
        1658 => "1111011011",  -- -1.1700
        1659 => "0000000001",  -- +0.0172
        1660 => "0000000111",  -- +0.2150
        1661 => "1111100000",  -- -1.0004
        1662 => "0000011010",  -- +0.8086
        1663 => "0000011100",  -- +0.8651
        1664 => "0000001010",  -- +0.2998
        1665 => "0000101011",  -- +1.3456
        1666 => "0000101000",  -- +1.2608
        1667 => "0000100001",  -- +1.0347
        1668 => "0000101000",  -- +1.2608
        1669 => "0000100101",  -- +1.1478
        1670 => "0000011001",  -- +0.7803
        1671 => "0000011101",  -- +0.8934
        1672 => "0000010110",  -- +0.6955
        1673 => "0000000111",  -- +0.2150
        1674 => "0000010100",  -- +0.6107
        1675 => "1111111001",  -- -0.2090
        1676 => "1111110111",  -- -0.2938
        1677 => "0000001111",  -- +0.4694
        1678 => "1111101001",  -- -0.7177
        1679 => "1111101011",  -- -0.6612
        1680 => "0000100000",  -- +1.0064
        1681 => "0000000010",  -- +0.0737
        1682 => "1111111101",  -- -0.0959
        1683 => "0000010000",  -- +0.4977
        1684 => "0000000001",  -- +0.0172
        1685 => "1111110010",  -- -0.4351
        1686 => "0000000101",  -- +0.1585
        1687 => "1111110101",  -- -0.3503
        1688 => "1111100011",  -- -0.9156
        1689 => "0000000100",  -- +0.1302
        1690 => "1111101111",  -- -0.5199
        1691 => "1111011111",  -- -1.0286
        1692 => "1111111100",  -- -0.1242
        1693 => "1111101000",  -- -0.7460
        1694 => "1111011001",  -- -1.2265
        1695 => "1111110101",  -- -0.3503
        1696 => "1111100001",  -- -0.9721
        1697 => "1111010010",  -- -1.4526
        1698 => "1111101110",  -- -0.5764
        1699 => "1111011011",  -- -1.1417
        1700 => "1111001101",  -- -1.5939
        1701 => "1111010011",  -- -1.3961
        1702 => "1111000011",  -- -1.9049
        1703 => "1110110101",  -- -2.3571
        1704 => "1111011111",  -- -1.0286
        1705 => "1111001111",  -- -1.5374
        1706 => "1111000000",  -- -1.9897
        1707 => "1111101110",  -- -0.5481
        1708 => "1111011111",  -- -1.0286
        1709 => "1111010001",  -- -1.4809
        1710 => "1111101100",  -- -0.6329
        1711 => "1111011100",  -- -1.1134
        1712 => "1111001111",  -- -1.5374
        1713 => "1111101000",  -- -0.7460
        1714 => "1111011000",  -- -1.2548
        1715 => "1111001011",  -- -1.6505
        1716 => "1111101011",  -- -0.6612
        1717 => "1111011011",  -- -1.1700
        1718 => "1111010000",  -- -1.5092
        1719 => "1111100000",  -- -1.0004
        1720 => "1111010000",  -- -1.5092
        1721 => "1111000101",  -- -1.8483
        1722 => "1111011011",  -- -1.1417
        1723 => "1111001010",  -- -1.6787
        1724 => "1110111111",  -- -2.0462
        1725 => "1111100001",  -- -0.9721
        1726 => "1111010000",  -- -1.5092
        1727 => "1111000011"   -- -1.9049
    );
    
begin
    
    process(clk)
    begin
        if rising_edge(clk) then
            dout_reg <= mem(to_integer(unsigned(addr)));
        end if;
    end process;

    -- Output assignment
    dout <= dout_reg;
end architecture rtl;
