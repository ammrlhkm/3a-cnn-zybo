--------------------------------------------------------------------------------
-- VHDL ROM with NORMALIZED image pixels (fixed-point format)
-- Generated from: 6_green_frog_s_000634.ppm
-- Generated on: 2025-12-18 08:57:09
-- 
-- Image size: 24x24 RGB
-- Memory depth: 1728 values
-- Address bits: 11
--
-- Normalization applied (matches cnn_ref.py):
--   mean = 90.2407
--   std_dev = 40.4184
--   normalized = (pixel - mean) / std_dev
--
-- Fixed-point format: Q5.5 (signed)
--   Total bits: 10
--   Integer bits: 5 (including sign)
--   Fractional bits: 5
--   Range: [-16.0000, 15.9688]
--   Resolution: 0.031250
--
-- Memory layout: Interleaved RGB
--   addr = (h * 24 + w) * 3 + channel
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity cnn_input_rom is
    generic (
        CELL_COUNT : integer := 1728;
        ADDR_WIDTH : integer := 11;
        DATA_WIDTH : integer := 10
    );
    port (
        clk     : in  std_logic;
        addr    : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        re      : in  std_logic;
        dout    : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end entity cnn_input_rom;

architecture rtl of cnn_input_rom is
    
    type mem_type is array (0 to CELL_COUNT-1) of std_logic_vector(DATA_WIDTH-1 downto 0);

    -- Output register for better timing (addresses SYNTH-6 warning)
    signal dout_reg : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');

    -- Normalized fixed-point pixel values
    constant mem : mem_type := (
        0 => "1111110011",  -- -0.4018
        1 => "1111111010",  -- -0.1791
        2 => "1111110001",  -- -0.4513
        3 => "1111111010",  -- -0.1791
        4 => "1111111111",  -- -0.0307
        5 => "1111110100",  -- -0.3523
        6 => "1111110100",  -- -0.3523
        7 => "1111111001",  -- -0.2039
        8 => "1111101111",  -- -0.5008
        9 => "1111100100",  -- -0.8719
        10 => "1111101001",  -- -0.6987
        11 => "1111011011",  -- -1.1441
        12 => "1111111010",  -- -0.1791
        13 => "0000000001",  -- +0.0435
        14 => "1111101000",  -- -0.7235
        15 => "1111111011",  -- -0.1544
        16 => "0000000011",  -- +0.1177
        17 => "1111100000",  -- -0.9709
        18 => "1111110011",  -- -0.3771
        19 => "1111111110",  -- -0.0554
        20 => "1111010011",  -- -1.3915
        21 => "1111110011",  -- -0.3771
        22 => "1111111110",  -- -0.0554
        23 => "1111001111",  -- -1.5152
        24 => "1111110110",  -- -0.3029
        25 => "0000000001",  -- +0.0435
        26 => "1111010001",  -- -1.4657
        27 => "1111111111",  -- -0.0307
        28 => "0000001010",  -- +0.3404
        29 => "1111010111",  -- -1.2678
        30 => "1111111111",  -- -0.0060
        31 => "0000001011",  -- +0.3652
        32 => "1111010110",  -- -1.2925
        33 => "1111111101",  -- -0.0802
        34 => "0000000111",  -- +0.2415
        35 => "1111010100",  -- -1.3667
        36 => "1111111010",  -- -0.1791
        37 => "0000000000",  -- +0.0188
        38 => "1111011001",  -- -1.2183
        39 => "1111101100",  -- -0.5997
        40 => "1111101111",  -- -0.5008
        41 => "1111011010",  -- -1.1688
        42 => "1111101101",  -- -0.5750
        43 => "1111101111",  -- -0.5255
        44 => "1111100101",  -- -0.8224
        45 => "1111101111",  -- -0.5008
        46 => "1111110001",  -- -0.4513
        47 => "1111100111",  -- -0.7729
        48 => "1111110110",  -- -0.3029
        49 => "1111110111",  -- -0.2534
        50 => "1111101000",  -- -0.7235
        51 => "1111110111",  -- -0.2534
        52 => "1111110101",  -- -0.3276
        53 => "1111101000",  -- -0.7235
        54 => "1111111011",  -- -0.1544
        55 => "1111110111",  -- -0.2534
        56 => "1111101100",  -- -0.6245
        57 => "1111111101",  -- -0.0802
        58 => "1111111010",  -- -0.1791
        59 => "1111101110",  -- -0.5503
        60 => "1111111101",  -- -0.0802
        61 => "1111111010",  -- -0.1791
        62 => "1111101110",  -- -0.5503
        63 => "1111111100",  -- -0.1049
        64 => "1111111000",  -- -0.2286
        65 => "1111101100",  -- -0.5997
        66 => "1111111111",  -- -0.0307
        67 => "1111111000",  -- -0.2286
        68 => "1111110000",  -- -0.4760
        69 => "1111111111",  -- -0.0307
        70 => "1111110111",  -- -0.2534
        71 => "1111110001",  -- -0.4513
        72 => "1111110010",  -- -0.4266
        73 => "1111111001",  -- -0.2039
        74 => "1111110000",  -- -0.4760
        75 => "1111110010",  -- -0.4266
        76 => "1111110111",  -- -0.2781
        77 => "1111101100",  -- -0.5997
        78 => "1111101111",  -- -0.5008
        79 => "1111110100",  -- -0.3523
        80 => "1111101001",  -- -0.6987
        81 => "1111101111",  -- -0.5008
        82 => "1111110101",  -- -0.3276
        83 => "1111100100",  -- -0.8472
        84 => "1111101111",  -- -0.5008
        85 => "1111110111",  -- -0.2534
        86 => "1111011011",  -- -1.1441
        87 => "1111101111",  -- -0.5255
        88 => "1111111001",  -- -0.2039
        89 => "1111010010",  -- -1.4162
        90 => "1111110000",  -- -0.4760
        91 => "1111111011",  -- -0.1297
        92 => "1111001101",  -- -1.5894
        93 => "1111110010",  -- -0.4266
        94 => "1111111101",  -- -0.0802
        95 => "1111001010",  -- -1.6636
        96 => "1111110011",  -- -0.3771
        97 => "1111111111",  -- -0.0060
        98 => "1111001001",  -- -1.6884
        99 => "1111110110",  -- -0.3029
        100 => "0000000010",  -- +0.0930
        101 => "1111001000",  -- -1.7378
        102 => "1111110110",  -- -0.3029
        103 => "0000000010",  -- +0.0930
        104 => "1111000100",  -- -1.8615
        105 => "1111111000",  -- -0.2286
        106 => "0000000011",  -- +0.1177
        107 => "1111000011",  -- -1.8863
        108 => "1111111111",  -- -0.0060
        109 => "0000000110",  -- +0.2167
        110 => "1111010001",  -- -1.4657
        111 => "1111111111",  -- -0.0307
        112 => "0000000010",  -- +0.0930
        113 => "1111100010",  -- -0.9214
        114 => "0000000100",  -- +0.1425
        115 => "0000000110",  -- +0.1920
        116 => "1111110111",  -- -0.2781
        117 => "0000000110",  -- +0.1920
        118 => "0000000110",  -- +0.2167
        119 => "1111111011",  -- -0.1544
        120 => "0000000111",  -- +0.2415
        121 => "0000000111",  -- +0.2415
        122 => "1111111010",  -- -0.1791
        123 => "0000001010",  -- +0.3404
        124 => "0000000111",  -- +0.2415
        125 => "1111111001",  -- -0.2039
        126 => "0000001001",  -- +0.2909
        127 => "0000000100",  -- +0.1425
        128 => "1111110110",  -- -0.3029
        129 => "0000001010",  -- +0.3404
        130 => "0000000110",  -- +0.1920
        131 => "1111110111",  -- -0.2534
        132 => "0000000110",  -- +0.2167
        133 => "0000000010",  -- +0.0683
        134 => "1111110100",  -- -0.3523
        135 => "0000000011",  -- +0.1177
        136 => "1111111110",  -- -0.0554
        137 => "1111110001",  -- -0.4513
        138 => "0000000101",  -- +0.1672
        139 => "1111111110",  -- -0.0554
        140 => "1111110101",  -- -0.3276
        141 => "0000000010",  -- +0.0930
        142 => "1111111010",  -- -0.1791
        143 => "1111110011",  -- -0.3771
        144 => "1111110011",  -- -0.4018
        145 => "1111111000",  -- -0.2286
        146 => "1111110000",  -- -0.4760
        147 => "1111101001",  -- -0.6987
        148 => "1111101000",  -- -0.7235
        149 => "1111100100",  -- -0.8719
        150 => "1111011010",  -- -1.1688
        151 => "1111011001",  -- -1.1935
        152 => "1111010001",  -- -1.4409
        153 => "1111100000",  -- -0.9709
        154 => "1111100100",  -- -0.8719
        155 => "1111010001",  -- -1.4409
        156 => "1111101110",  -- -0.5503
        157 => "1111111010",  -- -0.1791
        158 => "1111010110",  -- -1.2925
        159 => "1111101011",  -- -0.6492
        160 => "1111111101",  -- -0.0802
        161 => "1111001011",  -- -1.6389
        162 => "1111101110",  -- -0.5503
        163 => "1111111110",  -- -0.0554
        164 => "1111001000",  -- -1.7378
        165 => "1111110000",  -- -0.4760
        166 => "1111111111",  -- -0.0307
        167 => "1111000111",  -- -1.7626
        168 => "1111110011",  -- -0.3771
        169 => "0000000000",  -- +0.0188
        170 => "1111000110",  -- -1.7873
        171 => "1111110011",  -- -0.4018
        172 => "1111111101",  -- -0.0802
        173 => "1111000001",  -- -1.9605
        174 => "1111111000",  -- -0.2286
        175 => "0000000010",  -- +0.0683
        176 => "1111000011",  -- -1.8863
        177 => "0000000010",  -- +0.0930
        178 => "0000001000",  -- +0.2662
        179 => "1111001001",  -- -1.7131
        180 => "0000000100",  -- +0.1425
        181 => "0000000110",  -- +0.1920
        182 => "1111001011",  -- -1.6389
        183 => "0000000110",  -- +0.1920
        184 => "0000000111",  -- +0.2415
        185 => "1111011001",  -- -1.2183
        186 => "0000001111",  -- +0.4889
        187 => "0000010001",  -- +0.5384
        188 => "1111101111",  -- -0.5008
        189 => "0000010010",  -- +0.5878
        190 => "0000010011",  -- +0.6126
        191 => "1111111111",  -- -0.0307
        192 => "0000001001",  -- +0.2909
        193 => "0000001011",  -- +0.3652
        194 => "1111111100",  -- -0.1049
        195 => "0000000111",  -- +0.2415
        196 => "0000001010",  -- +0.3157
        197 => "1111110111",  -- -0.2534
        198 => "0000001010",  -- +0.3404
        199 => "0000001010",  -- +0.3157
        200 => "1111110111",  -- -0.2781
        201 => "0000001110",  -- +0.4641
        202 => "0000001010",  -- +0.3157
        203 => "1111111001",  -- -0.2039
        204 => "0000000110",  -- +0.2167
        205 => "0000000000",  -- +0.0188
        206 => "1111110011",  -- -0.3771
        207 => "0000000000",  -- +0.0188
        208 => "1111110111",  -- -0.2534
        209 => "1111110001",  -- -0.4513
        210 => "1111111011",  -- -0.1297
        211 => "1111110110",  -- -0.3029
        212 => "1111110001",  -- -0.4513
        213 => "1111110111",  -- -0.2534
        214 => "1111110011",  -- -0.4018
        215 => "1111101101",  -- -0.5750
        216 => "1111110000",  -- -0.4760
        217 => "1111110100",  -- -0.3523
        218 => "1111101101",  -- -0.5750
        219 => "1111100110",  -- -0.7977
        220 => "1111100100",  -- -0.8719
        221 => "1111100000",  -- -0.9709
        222 => "1111011001",  -- -1.1935
        223 => "1111010110",  -- -1.2925
        224 => "1111001110",  -- -1.5399
        225 => "1111011001",  -- -1.2183
        226 => "1111011011",  -- -1.1441
        227 => "1111000110",  -- -1.8121
        228 => "1111100101",  -- -0.8224
        229 => "1111110100",  -- -0.3523
        230 => "1111001010",  -- -1.6636
        231 => "1111100011",  -- -0.8966
        232 => "1111111011",  -- -0.1297
        233 => "1111000010",  -- -1.9358
        234 => "1111100110",  -- -0.7977
        235 => "1111111001",  -- -0.2039
        236 => "1111000000",  -- -1.9853
        237 => "1111101010",  -- -0.6740
        238 => "1111111000",  -- -0.2286
        239 => "1111000001",  -- -1.9605
        240 => "1111101100",  -- -0.6245
        241 => "1111110111",  -- -0.2534
        242 => "1110111111",  -- -2.0100
        243 => "1111110000",  -- -0.4760
        244 => "1111111010",  -- -0.1791
        245 => "1111000001",  -- -1.9605
        246 => "1111111001",  -- -0.2039
        247 => "0000000000",  -- +0.0188
        248 => "1111000110",  -- -1.8121
        249 => "0000000100",  -- +0.1425
        250 => "0000000110",  -- +0.2167
        251 => "1111001011",  -- -1.6389
        252 => "0000001011",  -- +0.3652
        253 => "0000001010",  -- +0.3157
        254 => "1111001110",  -- -1.5399
        255 => "0000000010",  -- +0.0930
        256 => "0000000100",  -- +0.1425
        257 => "1111001001",  -- -1.6884
        258 => "0000000010",  -- +0.0683
        259 => "0000000101",  -- +0.1672
        260 => "1111010010",  -- -1.4162
        261 => "0000001010",  -- +0.3157
        262 => "0000001110",  -- +0.4394
        263 => "1111101010",  -- -0.6740
        264 => "0000001010",  -- +0.3157
        265 => "0000001110",  -- +0.4641
        266 => "1111110101",  -- -0.3276
        267 => "0000001100",  -- +0.3899
        268 => "0000010010",  -- +0.5878
        269 => "1111110111",  -- -0.2781
        270 => "0000001110",  -- +0.4394
        271 => "0000010010",  -- +0.5631
        272 => "1111110101",  -- -0.3276
        273 => "0000000101",  -- +0.1672
        274 => "0000000010",  -- +0.0930
        275 => "1111101011",  -- -0.6492
        276 => "0000000010",  -- +0.0683
        277 => "1111111001",  -- -0.2039
        278 => "1111101100",  -- -0.6245
        279 => "0000000000",  -- +0.0188
        280 => "1111110101",  -- -0.3276
        281 => "1111110010",  -- -0.4266
        282 => "1111111011",  -- -0.1544
        283 => "1111110101",  -- -0.3276
        284 => "1111110001",  -- -0.4513
        285 => "1111110111",  -- -0.2534
        286 => "1111110011",  -- -0.3771
        287 => "1111101100",  -- -0.5997
        288 => "1111111110",  -- -0.0554
        289 => "0000000010",  -- +0.0930
        290 => "1111111001",  -- -0.2039
        291 => "0000001010",  -- +0.3157
        292 => "0000001010",  -- +0.3404
        293 => "0000000010",  -- +0.0683
        294 => "1111111101",  -- -0.0802
        295 => "1111111011",  -- -0.1297
        296 => "1111101111",  -- -0.5008
        297 => "1111011100",  -- -1.0946
        298 => "1111011111",  -- -1.0203
        299 => "1111000111",  -- -1.7626
        300 => "1111100100",  -- -0.8472
        301 => "1111110010",  -- -0.4266
        302 => "1111000110",  -- -1.7873
        303 => "1111100100",  -- -0.8472
        304 => "1111111011",  -- -0.1544
        305 => "1111000010",  -- -1.9358
        306 => "1111101111",  -- -0.5255
        307 => "0000000000",  -- +0.0188
        308 => "1111001100",  -- -1.6141
        309 => "1111111001",  -- -0.2039
        310 => "0000000110",  -- +0.2167
        311 => "1111010101",  -- -1.3172
        312 => "1111111000",  -- -0.2286
        313 => "0000000101",  -- +0.1672
        314 => "1111010001",  -- -1.4409
        315 => "1111111101",  -- -0.0802
        316 => "0000000111",  -- +0.2415
        317 => "1111010010",  -- -1.4162
        318 => "1111111111",  -- -0.0060
        319 => "0000001000",  -- +0.2662
        320 => "1111010010",  -- -1.4162
        321 => "1111111101",  -- -0.0802
        322 => "0000000010",  -- +0.0930
        323 => "1111001000",  -- -1.7378
        324 => "0000000110",  -- +0.1920
        325 => "0000001000",  -- +0.2662
        326 => "1111001001",  -- -1.6884
        327 => "0000000110",  -- +0.2167
        328 => "0000001010",  -- +0.3404
        329 => "1111001011",  -- -1.6389
        330 => "0000000010",  -- +0.0930
        331 => "0000001000",  -- +0.2662
        332 => "1111001100",  -- -1.6141
        333 => "0000000000",  -- +0.0188
        334 => "0000000110",  -- +0.1920
        335 => "1111010010",  -- -1.4162
        336 => "0000000101",  -- +0.1672
        337 => "0000001100",  -- +0.3899
        338 => "1111011111",  -- -1.0203
        339 => "0000001001",  -- +0.2909
        340 => "0000010000",  -- +0.5136
        341 => "1111100100",  -- -0.8472
        342 => "0000001100",  -- +0.3899
        343 => "0000010010",  -- +0.5878
        344 => "1111101000",  -- -0.7482
        345 => "0000001001",  -- +0.2909
        346 => "0000001010",  -- +0.3157
        347 => "1111100111",  -- -0.7729
        348 => "0000000010",  -- +0.0930
        349 => "1111111101",  -- -0.0802
        350 => "1111100111",  -- -0.7729
        351 => "0000000110",  -- +0.2167
        352 => "1111111011",  -- -0.1297
        353 => "1111110011",  -- -0.3771
        354 => "0000000101",  -- +0.1672
        355 => "1111111001",  -- -0.2039
        356 => "1111110010",  -- -0.4266
        357 => "0000000001",  -- +0.0435
        358 => "1111110110",  -- -0.3029
        359 => "1111101010",  -- -0.6740
        360 => "0000100100",  -- +1.1321
        361 => "0000101000",  -- +1.2806
        362 => "0000011101",  -- +0.9342
        363 => "0000110001",  -- +1.5527
        364 => "0000110100",  -- +1.6517
        365 => "0000101000",  -- +1.2558
        366 => "0000001010",  -- +0.3404
        367 => "0000001010",  -- +0.3404
        368 => "1111111011",  -- -0.1297
        369 => "1111100000",  -- -0.9709
        370 => "1111100011",  -- -0.8966
        371 => "1111001001",  -- -1.6884
        372 => "1111101000",  -- -0.7482
        373 => "1111110011",  -- -0.3771
        374 => "1111001001",  -- -1.7131
        375 => "1111100111",  -- -0.7729
        376 => "1111111011",  -- -0.1544
        377 => "1111000100",  -- -1.8615
        378 => "1111110010",  -- -0.4266
        379 => "0000000010",  -- +0.0683
        380 => "1111010010",  -- -1.4162
        381 => "0000000101",  -- +0.1672
        382 => "0000010010",  -- +0.5631
        383 => "1111100100",  -- -0.8472
        384 => "0000001000",  -- +0.2662
        385 => "0000010101",  -- +0.6621
        386 => "1111100101",  -- -0.8224
        387 => "0000001110",  -- +0.4394
        388 => "0000011010",  -- +0.8352
        389 => "1111101000",  -- -0.7235
        390 => "0000001001",  -- +0.2909
        391 => "0000010101",  -- +0.6621
        392 => "1111100010",  -- -0.9214
        393 => "1111111111",  -- -0.0060
        394 => "0000001000",  -- +0.2662
        395 => "1111001110",  -- -1.5399
        396 => "0000000011",  -- +0.1177
        397 => "0000001010",  -- +0.3157
        398 => "1111001001",  -- -1.7131
        399 => "0000000101",  -- +0.1672
        400 => "0000001100",  -- +0.3899
        401 => "1111001001",  -- -1.6884
        402 => "0000000101",  -- +0.1672
        403 => "0000001101",  -- +0.4146
        404 => "1111001001",  -- -1.6884
        405 => "0000000010",  -- +0.0683
        406 => "0000001010",  -- +0.3157
        407 => "1111001000",  -- -1.7378
        408 => "0000000010",  -- +0.0683
        409 => "0000001010",  -- +0.3404
        410 => "1111001011",  -- -1.6389
        411 => "0000000110",  -- +0.2167
        412 => "0000001111",  -- +0.4889
        413 => "1111010100",  -- -1.3667
        414 => "0000001011",  -- +0.3652
        415 => "0000010100",  -- +0.6373
        416 => "1111011100",  -- -1.1193
        417 => "0000001111",  -- +0.4889
        418 => "0000010101",  -- +0.6868
        419 => "1111100110",  -- -0.7977
        420 => "0000001010",  -- +0.3157
        421 => "0000000111",  -- +0.2415
        422 => "1111101000",  -- -0.7235
        423 => "0000001011",  -- +0.3652
        424 => "1111111111",  -- -0.0060
        425 => "1111110001",  -- -0.4513
        426 => "0000001110",  -- +0.4394
        427 => "1111111011",  -- -0.1297
        428 => "1111101111",  -- -0.5008
        429 => "0000001110",  -- +0.4394
        430 => "1111111011",  -- -0.1544
        431 => "1111101100",  -- -0.6245
        432 => "0000110111",  -- +1.7259
        433 => "0000111011",  -- +1.8744
        434 => "0000110000",  -- +1.5280
        435 => "0000111000",  -- +1.7754
        436 => "0000111111",  -- +1.9733
        437 => "0000110000",  -- +1.5280
        438 => "1111111101",  -- -0.0802
        439 => "1111111111",  -- -0.0307
        440 => "1111110000",  -- -0.4760
        441 => "1111100000",  -- -0.9956
        442 => "1111100010",  -- -0.9214
        443 => "1111001011",  -- -1.6389
        444 => "1111101101",  -- -0.5750
        445 => "1111110111",  -- -0.2534
        446 => "1111010000",  -- -1.4904
        447 => "1111100100",  -- -0.8472
        448 => "1111110101",  -- -0.3276
        449 => "1111000110",  -- -1.8121
        450 => "1111100010",  -- -0.9214
        451 => "1111101111",  -- -0.5008
        452 => "1111001001",  -- -1.7131
        453 => "1111111110",  -- -0.0554
        454 => "0000001010",  -- +0.3404
        455 => "1111011111",  -- -1.0203
        456 => "0000001000",  -- +0.2662
        457 => "0000010110",  -- +0.7115
        458 => "1111101000",  -- -0.7482
        459 => "0000010001",  -- +0.5384
        460 => "0000011111",  -- +0.9837
        461 => "1111101110",  -- -0.5503
        462 => "0000001101",  -- +0.4146
        463 => "0000011101",  -- +0.9095
        464 => "1111101010",  -- -0.6740
        465 => "1111111111",  -- -0.0060
        466 => "0000001101",  -- +0.4146
        467 => "1111010010",  -- -1.4162
        468 => "0000000010",  -- +0.0930
        469 => "0000001100",  -- +0.3899
        470 => "1111001100",  -- -1.6141
        471 => "0000000100",  -- +0.1425
        472 => "0000001110",  -- +0.4394
        473 => "1111001101",  -- -1.5647
        474 => "0000000010",  -- +0.0930
        475 => "0000001011",  -- +0.3652
        476 => "1111001001",  -- -1.7131
        477 => "0000000100",  -- +0.1425
        478 => "0000001100",  -- +0.3899
        479 => "1111000110",  -- -1.8121
        480 => "0000000100",  -- +0.1425
        481 => "0000001100",  -- +0.3899
        482 => "1111000100",  -- -1.8615
        483 => "0000000011",  -- +0.1177
        484 => "0000001011",  -- +0.3652
        485 => "1111001000",  -- -1.7378
        486 => "0000000100",  -- +0.1425
        487 => "0000001111",  -- +0.4889
        488 => "1111001110",  -- -1.5399
        489 => "0000001000",  -- +0.2662
        490 => "0000010010",  -- +0.5878
        491 => "1111011010",  -- -1.1688
        492 => "0000001010",  -- +0.3404
        493 => "0000001011",  -- +0.3652
        494 => "1111100100",  -- -0.8719
        495 => "0000010010",  -- +0.5631
        496 => "0000000110",  -- +0.1920
        497 => "1111101111",  -- -0.5008
        498 => "0000011011",  -- +0.8600
        499 => "0000000110",  -- +0.1920
        500 => "1111110101",  -- -0.3276
        501 => "0000011100",  -- +0.8847
        502 => "0000000100",  -- +0.1425
        503 => "1111110011",  -- -0.4018
        504 => "0000110111",  -- +1.7259
        505 => "0000111100",  -- +1.8991
        506 => "0000110001",  -- +1.5527
        507 => "0000110110",  -- +1.7012
        508 => "0000111110",  -- +1.9486
        509 => "0000110001",  -- +1.5527
        510 => "1111111111",  -- -0.0060
        511 => "0000000010",  -- +0.0683
        512 => "1111110111",  -- -0.2781
        513 => "1111011011",  -- -1.1441
        514 => "1111011100",  -- -1.0946
        515 => "1111001010",  -- -1.6636
        516 => "1111110001",  -- -0.4513
        517 => "1111111000",  -- -0.2286
        518 => "1111011000",  -- -1.2430
        519 => "1111101111",  -- -0.5255
        520 => "1111111100",  -- -0.1049
        521 => "1111010011",  -- -1.3915
        522 => "1111100110",  -- -0.7977
        523 => "1111110011",  -- -0.4018
        524 => "1111001100",  -- -1.6141
        525 => "1111111100",  -- -0.1049
        526 => "0000001010",  -- +0.3157
        527 => "1111011100",  -- -1.0946
        528 => "0000001010",  -- +0.3157
        529 => "0000011001",  -- +0.8105
        530 => "1111101000",  -- -0.7235
        531 => "1111111111",  -- -0.0060
        532 => "0000010001",  -- +0.5384
        533 => "1111011110",  -- -1.0451
        534 => "0000000101",  -- +0.1672
        535 => "0000011001",  -- +0.7858
        536 => "1111100100",  -- -0.8719
        537 => "0000000001",  -- +0.0435
        538 => "0000010010",  -- +0.5878
        539 => "1111010111",  -- -1.2678
        540 => "1111111111",  -- -0.0060
        541 => "0000001100",  -- +0.3899
        542 => "1111001111",  -- -1.5152
        543 => "0000000100",  -- +0.1425
        544 => "0000001110",  -- +0.4641
        545 => "1111010101",  -- -1.3420
        546 => "0000000011",  -- +0.1177
        547 => "0000001100",  -- +0.3899
        548 => "1111010001",  -- -1.4657
        549 => "0000000010",  -- +0.0930
        550 => "0000001010",  -- +0.3157
        551 => "1111001001",  -- -1.7131
        552 => "0000000110",  -- +0.2167
        553 => "0000001101",  -- +0.4146
        554 => "1111000111",  -- -1.7626
        555 => "0000000110",  -- +0.1920
        556 => "0000001011",  -- +0.3652
        557 => "1111001001",  -- -1.7131
        558 => "1111111101",  -- -0.0802
        559 => "0000001010",  -- +0.3157
        560 => "1111000110",  -- -1.7873
        561 => "0000000001",  -- +0.0435
        562 => "0000001111",  -- +0.4889
        563 => "1111010001",  -- -1.4657
        564 => "0000000101",  -- +0.1672
        565 => "0000001001",  -- +0.2909
        566 => "1111011001",  -- -1.1935
        567 => "0000010001",  -- +0.5384
        568 => "0000000101",  -- +0.1672
        569 => "1111100111",  -- -0.7729
        570 => "0000100000",  -- +1.0084
        571 => "0000001000",  -- +0.2662
        572 => "1111110100",  -- -0.3523
        573 => "0000100000",  -- +1.0084
        574 => "0000000110",  -- +0.2167
        575 => "1111110101",  -- -0.3276
        576 => "0000110000",  -- +1.5280
        577 => "0000110101",  -- +1.6764
        578 => "0000101100",  -- +1.3796
        579 => "0000101101",  -- +1.4290
        580 => "0000110110",  -- +1.7012
        581 => "0000101100",  -- +1.3796
        582 => "0000010010",  -- +0.5878
        583 => "0000010101",  -- +0.6621
        584 => "0000001101",  -- +0.4146
        585 => "1111011110",  -- -1.0451
        586 => "1111011110",  -- -1.0451
        587 => "1111010001",  -- -1.4409
        588 => "1111101110",  -- -0.5503
        589 => "1111110010",  -- -0.4266
        590 => "1111011010",  -- -1.1688
        591 => "1111111110",  -- -0.0554
        592 => "0000001000",  -- +0.2662
        593 => "1111100100",  -- -0.8719
        594 => "0000000010",  -- +0.0930
        595 => "0000001110",  -- +0.4394
        596 => "1111100001",  -- -0.9461
        597 => "0000001010",  -- +0.3157
        598 => "0000010111",  -- +0.7363
        599 => "1111100111",  -- -0.7729
        600 => "0000010011",  -- +0.6126
        601 => "0000100011",  -- +1.1074
        602 => "1111110000",  -- -0.4760
        603 => "0000000100",  -- +0.1425
        604 => "0000010111",  -- +0.7363
        605 => "1111100001",  -- -0.9461
        606 => "1111111110",  -- -0.0554
        607 => "0000010100",  -- +0.6373
        608 => "1111011011",  -- -1.1441
        609 => "0000000010",  -- +0.0683
        610 => "0000010101",  -- +0.6621
        611 => "1111011001",  -- -1.2183
        612 => "1111111111",  -- -0.0307
        613 => "0000001101",  -- +0.4146
        614 => "1111010011",  -- -1.3915
        615 => "0000001000",  -- +0.2662
        616 => "0000010011",  -- +0.6126
        617 => "1111100000",  -- -0.9956
        618 => "0000000110",  -- +0.1920
        619 => "0000001110",  -- +0.4394
        620 => "1111011011",  -- -1.1441
        621 => "0000000010",  -- +0.0930
        622 => "0000001001",  -- +0.2909
        623 => "1111010000",  -- -1.4904
        624 => "0000000110",  -- +0.2167
        625 => "0000001011",  -- +0.3652
        626 => "1111001101",  -- -1.5894
        627 => "0000001000",  -- +0.2662
        628 => "0000001100",  -- +0.3899
        629 => "1111001110",  -- -1.5399
        630 => "1111111011",  -- -0.1544
        631 => "0000000111",  -- +0.2415
        632 => "1111000110",  -- -1.7873
        633 => "1111111011",  -- -0.1297
        634 => "0000001011",  -- +0.3652
        635 => "1111001100",  -- -1.6141
        636 => "0000001011",  -- +0.3652
        637 => "0000010001",  -- +0.5384
        638 => "1111011100",  -- -1.0946
        639 => "0000001111",  -- +0.4889
        640 => "0000000100",  -- +0.1425
        641 => "1111100000",  -- -0.9956
        642 => "0000011011",  -- +0.8600
        643 => "0000000100",  -- +0.1425
        644 => "1111101111",  -- -0.5255
        645 => "0000100001",  -- +1.0332
        646 => "0000001000",  -- +0.2662
        647 => "1111111000",  -- -0.2286
        648 => "0000101010",  -- +1.3301
        649 => "0000101100",  -- +1.4043
        650 => "0000100101",  -- +1.1816
        651 => "0000101000",  -- +1.2806
        652 => "0000101100",  -- +1.4043
        653 => "0000100101",  -- +1.1569
        654 => "0000100100",  -- +1.1321
        655 => "0000100011",  -- +1.1074
        656 => "0000011100",  -- +0.8847
        657 => "1111110111",  -- -0.2534
        658 => "1111110100",  -- -0.3523
        659 => "1111101011",  -- -0.6492
        660 => "1111011101",  -- -1.0698
        661 => "1111011011",  -- -1.1441
        662 => "1111001101",  -- -1.5894
        663 => "1111110001",  -- -0.4513
        664 => "1111110010",  -- -0.4266
        665 => "1111011100",  -- -1.0946
        666 => "0000000010",  -- +0.0930
        667 => "0000001010",  -- +0.3157
        668 => "1111101000",  -- -0.7235
        669 => "0000001010",  -- +0.3404
        670 => "0000010101",  -- +0.6621
        671 => "1111101100",  -- -0.6245
        672 => "0000010010",  -- +0.5878
        673 => "0000100000",  -- +1.0084
        674 => "1111101111",  -- -0.5008
        675 => "0000010010",  -- +0.5631
        676 => "0000100001",  -- +1.0579
        677 => "1111101011",  -- -0.6492
        678 => "0000000001",  -- +0.0435
        679 => "0000010011",  -- +0.6126
        680 => "1111011000",  -- -1.2430
        681 => "0000000010",  -- +0.0930
        682 => "0000010010",  -- +0.5631
        683 => "1111010101",  -- -1.3420
        684 => "0000000010",  -- +0.0683
        685 => "0000001110",  -- +0.4394
        686 => "1111010101",  -- -1.3420
        687 => "0000001010",  -- +0.3157
        688 => "0000010110",  -- +0.7115
        689 => "1111100011",  -- -0.8966
        690 => "0000000101",  -- +0.1672
        691 => "0000010010",  -- +0.5631
        692 => "1111100000",  -- -0.9709
        693 => "0000000010",  -- +0.0683
        694 => "0000001101",  -- +0.4146
        695 => "1111011000",  -- -1.2430
        696 => "0000000100",  -- +0.1425
        697 => "0000001100",  -- +0.3899
        698 => "1111010010",  -- -1.4162
        699 => "0000000101",  -- +0.1672
        700 => "0000001100",  -- +0.3899
        701 => "1111001111",  -- -1.5152
        702 => "1111111011",  -- -0.1297
        703 => "0000001000",  -- +0.2662
        704 => "1111000110",  -- -1.7873
        705 => "1111111001",  -- -0.2039
        706 => "0000000111",  -- +0.2415
        707 => "1111000111",  -- -1.7626
        708 => "0000001101",  -- +0.4146
        709 => "0000010101",  -- +0.6621
        710 => "1111011101",  -- -1.0698
        711 => "0000001101",  -- +0.4146
        712 => "0000001011",  -- +0.3652
        713 => "1111100000",  -- -0.9709
        714 => "0000010000",  -- +0.5136
        715 => "0000000010",  -- +0.0683
        716 => "1111101000",  -- -0.7482
        717 => "0000011000",  -- +0.7610
        718 => "0000000110",  -- +0.1920
        719 => "1111110110",  -- -0.3029
        720 => "0000101000",  -- +1.2806
        721 => "0000101001",  -- +1.3053
        722 => "0000100010",  -- +1.0827
        723 => "0000101100",  -- +1.4043
        724 => "0000101101",  -- +1.4290
        725 => "0000100100",  -- +1.1321
        726 => "0000110000",  -- +1.5033
        727 => "0000101110",  -- +1.4538
        728 => "0000100101",  -- +1.1569
        729 => "0000100101",  -- +1.1569
        730 => "0000100000",  -- +1.0084
        731 => "0000010110",  -- +0.7115
        732 => "0000000010",  -- +0.0683
        733 => "1111111011",  -- -0.1544
        734 => "1111110000",  -- -0.4760
        735 => "1111110010",  -- -0.4266
        736 => "1111101100",  -- -0.6245
        737 => "1111011111",  -- -1.0203
        738 => "1111100000",  -- -0.9956
        739 => "1111100010",  -- -0.9214
        740 => "1111001101",  -- -1.5647
        741 => "1111101001",  -- -0.6987
        742 => "1111101111",  -- -0.5008
        743 => "1111010010",  -- -1.4162
        744 => "1111111111",  -- -0.0307
        745 => "0000000110",  -- +0.2167
        746 => "1111011100",  -- -1.0946
        747 => "0000000010",  -- +0.0930
        748 => "0000001101",  -- +0.4146
        749 => "1111011001",  -- -1.1935
        750 => "1111111111",  -- -0.0060
        751 => "0000001010",  -- +0.3404
        752 => "1111010001",  -- -1.4409
        753 => "0000000110",  -- +0.1920
        754 => "0000001110",  -- +0.4641
        755 => "1111010011",  -- -1.3915
        756 => "0000001001",  -- +0.2909
        757 => "0000010010",  -- +0.5878
        758 => "1111011000",  -- -1.2430
        759 => "0000001011",  -- +0.3652
        760 => "0000011010",  -- +0.8352
        761 => "1111100101",  -- -0.8224
        762 => "0000001010",  -- +0.3157
        763 => "0000011011",  -- +0.8600
        764 => "1111101000",  -- -0.7235
        765 => "0000000101",  -- +0.1672
        766 => "0000010101",  -- +0.6621
        767 => "1111100000",  -- -0.9956
        768 => "0000000010",  -- +0.0930
        769 => "0000001111",  -- +0.4889
        770 => "1111010111",  -- -1.2678
        771 => "0000000010",  -- +0.0930
        772 => "0000001110",  -- +0.4394
        773 => "1111001110",  -- -1.5399
        774 => "1111111100",  -- -0.1049
        775 => "0000001000",  -- +0.2662
        776 => "1111000110",  -- -1.8121
        777 => "1111111010",  -- -0.1791
        778 => "0000000110",  -- +0.1920
        779 => "1111000110",  -- -1.8121
        780 => "0000000011",  -- +0.1177
        781 => "0000001110",  -- +0.4394
        782 => "1111010101",  -- -1.3420
        783 => "0000001000",  -- +0.2662
        784 => "0000010000",  -- +0.5136
        785 => "1111100000",  -- -0.9709
        786 => "0000000001",  -- +0.0435
        787 => "1111111110",  -- -0.0554
        788 => "1111011110",  -- -1.0451
        789 => "0000001001",  -- +0.2909
        790 => "1111111111",  -- -0.0060
        791 => "1111101100",  -- -0.6245
        792 => "0000110000",  -- +1.5280
        793 => "0000110001",  -- +1.5527
        794 => "0000100111",  -- +1.2311
        795 => "0000110110",  -- +1.7012
        796 => "0000110111",  -- +1.7259
        797 => "0000101011",  -- +1.3548
        798 => "0000110010",  -- +1.5775
        799 => "0000110001",  -- +1.5527
        800 => "0000100100",  -- +1.1321
        801 => "0000110000",  -- +1.5280
        802 => "0000101100",  -- +1.4043
        803 => "0000011110",  -- +0.9590
        804 => "0000110101",  -- +1.6764
        805 => "0000110000",  -- +1.5033
        806 => "0000100001",  -- +1.0332
        807 => "0000010101",  -- +0.6868
        808 => "0000010000",  -- +0.5136
        809 => "1111111111",  -- -0.0060
        810 => "1111100010",  -- -0.9214
        811 => "1111100001",  -- -0.9461
        812 => "1111010000",  -- -1.4904
        813 => "1111100101",  -- -0.8224
        814 => "1111100110",  -- -0.7977
        815 => "1111010000",  -- -1.4904
        816 => "0000001010",  -- +0.3157
        817 => "0000001100",  -- +0.3899
        818 => "1111101011",  -- -0.6492
        819 => "0000000111",  -- +0.2415
        820 => "0000001010",  -- +0.3404
        821 => "1111100000",  -- -0.9709
        822 => "0000000011",  -- +0.1177
        823 => "0000001000",  -- +0.2662
        824 => "1111010111",  -- -1.2678
        825 => "0000001001",  -- +0.2909
        826 => "0000001111",  -- +0.4889
        827 => "1111010111",  -- -1.2678
        828 => "0000001111",  -- +0.4889
        829 => "0000011001",  -- +0.8105
        830 => "1111011111",  -- -1.0203
        831 => "0000010100",  -- +0.6373
        832 => "0000100101",  -- +1.1569
        833 => "1111101111",  -- -0.5255
        834 => "0000010000",  -- +0.5136
        835 => "0000100011",  -- +1.1074
        836 => "1111101111",  -- -0.5255
        837 => "0000001100",  -- +0.3899
        838 => "0000011101",  -- +0.9342
        839 => "1111101000",  -- -0.7235
        840 => "0000000101",  -- +0.1672
        841 => "0000010011",  -- +0.6126
        842 => "1111011011",  -- -1.1441
        843 => "0000000000",  -- +0.0188
        844 => "0000001110",  -- +0.4394
        845 => "1111001110",  -- -1.5399
        846 => "1111111101",  -- -0.0802
        847 => "0000001010",  -- +0.3404
        848 => "1111001000",  -- -1.7378
        849 => "1111111011",  -- -0.1297
        850 => "0000001000",  -- +0.2662
        851 => "1111000111",  -- -1.7626
        852 => "1111111011",  -- -0.1544
        853 => "0000000110",  -- +0.2167
        854 => "1111001100",  -- -1.6141
        855 => "0000000110",  -- +0.1920
        856 => "0000010000",  -- +0.5136
        857 => "1111011110",  -- -1.0451
        858 => "1111111011",  -- -0.1297
        859 => "1111111111",  -- -0.0307
        860 => "1111011001",  -- -1.2183
        861 => "1111111010",  -- -0.1791
        862 => "1111110110",  -- -0.3029
        863 => "1111011100",  -- -1.1193
        864 => "0000111010",  -- +1.8249
        865 => "0000111010",  -- +1.8249
        866 => "0000101110",  -- +1.4538
        867 => "0000111000",  -- +1.7507
        868 => "0000110111",  -- +1.7259
        869 => "0000101011",  -- +1.3548
        870 => "0000100101",  -- +1.1569
        871 => "0000100100",  -- +1.1321
        872 => "0000010101",  -- +0.6621
        873 => "0000010011",  -- +0.6126
        874 => "0000010010",  -- +0.5878
        875 => "1111111111",  -- -0.0060
        876 => "0000110100",  -- +1.6517
        877 => "0000110011",  -- +1.6022
        878 => "0000011101",  -- +0.9342
        879 => "0000101011",  -- +1.3548
        880 => "0000101001",  -- +1.3053
        881 => "0000010010",  -- +0.5878
        882 => "0000011101",  -- +0.9342
        883 => "0000011001",  -- +0.7858
        884 => "0000000110",  -- +0.1920
        885 => "0000001111",  -- +0.4889
        886 => "0000001010",  -- +0.3404
        887 => "1111110111",  -- -0.2534
        888 => "0000011001",  -- +0.8105
        889 => "0000010101",  -- +0.6868
        890 => "1111111101",  -- -0.0802
        891 => "0000011001",  -- +0.7858
        892 => "0000010110",  -- +0.7115
        893 => "1111110101",  -- -0.3276
        894 => "0000001010",  -- +0.3404
        895 => "0000001001",  -- +0.2909
        896 => "1111011111",  -- -1.0203
        897 => "0000001010",  -- +0.3157
        898 => "0000001110",  -- +0.4394
        899 => "1111011000",  -- -1.2430
        900 => "0000001011",  -- +0.3652
        901 => "0000010111",  -- +0.7363
        902 => "1111011100",  -- -1.0946
        903 => "0000001110",  -- +0.4641
        904 => "0000100001",  -- +1.0332
        905 => "1111101010",  -- -0.6740
        906 => "0000001110",  -- +0.4394
        907 => "0000100001",  -- +1.0579
        908 => "1111101110",  -- -0.5503
        909 => "0000001010",  -- +0.3404
        910 => "0000011101",  -- +0.9342
        911 => "1111101000",  -- -0.7482
        912 => "0000000101",  -- +0.1672
        913 => "0000010101",  -- +0.6621
        914 => "1111011100",  -- -1.1193
        915 => "1111111111",  -- -0.0060
        916 => "0000001110",  -- +0.4641
        917 => "1111010001",  -- -1.4657
        918 => "1111111110",  -- -0.0554
        919 => "0000001101",  -- +0.4146
        920 => "1111001100",  -- -1.6141
        921 => "1111111101",  -- -0.0802
        922 => "0000001100",  -- +0.3899
        923 => "1111001010",  -- -1.6636
        924 => "1111110111",  -- -0.2781
        925 => "0000000101",  -- +0.1672
        926 => "1111001001",  -- -1.7131
        927 => "0000000001",  -- +0.0435
        928 => "0000001110",  -- +0.4394
        929 => "1111011001",  -- -1.1935
        930 => "1111111101",  -- -0.0802
        931 => "0000000110",  -- +0.1920
        932 => "1111011010",  -- -1.1688
        933 => "1111111011",  -- -0.1297
        934 => "1111111100",  -- -0.1049
        935 => "1111011100",  -- -1.1193
        936 => "0000111111",  -- +1.9733
        937 => "0000111100",  -- +1.8991
        938 => "0000110010",  -- +1.5775
        939 => "0001000110",  -- +2.1960
        940 => "0001000100",  -- +2.1465
        941 => "0000111010",  -- +1.8249
        942 => "0001000011",  -- +2.1218
        943 => "0001000011",  -- +2.1218
        944 => "0000110101",  -- +1.6764
        945 => "0000011101",  -- +0.9095
        946 => "0000011110",  -- +0.9590
        947 => "0000001010",  -- +0.3404
        948 => "0001000011",  -- +2.1218
        949 => "0001000110",  -- +2.1960
        950 => "0000101110",  -- +1.4538
        951 => "0001010100",  -- +2.6414
        952 => "0001010110",  -- +2.6908
        953 => "0000111011",  -- +1.8744
        954 => "0000110100",  -- +1.6517
        955 => "0000110000",  -- +1.5033
        956 => "0000011001",  -- +0.7858
        957 => "0000110000",  -- +1.5280
        958 => "0000101000",  -- +1.2806
        959 => "0000010110",  -- +0.7115
        960 => "0000010010",  -- +0.5631
        961 => "0000001010",  -- +0.3404
        962 => "1111110111",  -- -0.2534
        963 => "0000101011",  -- +1.3548
        964 => "0000100101",  -- +1.1569
        965 => "0000001010",  -- +0.3157
        966 => "0000011101",  -- +0.9342
        967 => "0000011001",  -- +0.8105
        968 => "1111110011",  -- -0.3771
        969 => "0000001010",  -- +0.3157
        970 => "0000001110",  -- +0.4394
        971 => "1111011001",  -- -1.2183
        972 => "0000001010",  -- +0.3157
        973 => "0000011000",  -- +0.7610
        974 => "1111011100",  -- -1.1193
        975 => "0000001000",  -- +0.2662
        976 => "0000011100",  -- +0.8847
        977 => "1111100100",  -- -0.8472
        978 => "0000001010",  -- +0.3404
        979 => "0000100000",  -- +1.0084
        980 => "1111101100",  -- -0.6245
        981 => "0000001001",  -- +0.2909
        982 => "0000011101",  -- +0.9342
        983 => "1111101000",  -- -0.7482
        984 => "0000000101",  -- +0.1672
        985 => "0000010110",  -- +0.7115
        986 => "1111011110",  -- -1.0451
        987 => "0000000011",  -- +0.1177
        988 => "0000010011",  -- +0.6126
        989 => "1111011000",  -- -1.2430
        990 => "0000000000",  -- +0.0188
        991 => "0000010001",  -- +0.5384
        992 => "1111010001",  -- -1.4657
        993 => "1111111111",  -- -0.0307
        994 => "0000001111",  -- +0.4889
        995 => "1111001101",  -- -1.5647
        996 => "1111110111",  -- -0.2781
        997 => "0000000110",  -- +0.2167
        998 => "1111001001",  -- -1.7131
        999 => "1111111100",  -- -0.1049
        1000 => "0000001011",  -- +0.3652
        1001 => "1111010100",  -- -1.3667
        1002 => "0000000000",  -- +0.0188
        1003 => "0000001100",  -- +0.3899
        1004 => "1111011101",  -- -1.0698
        1005 => "0000000000",  -- +0.0188
        1006 => "0000000010",  -- +0.0930
        1007 => "1111100000",  -- -0.9956
        1008 => "0001100111",  -- +3.2351
        1009 => "0001100101",  -- +3.1609
        1010 => "0001011110",  -- +2.9630
        1011 => "0001110100",  -- +3.6557
        1012 => "0001110011",  -- +3.6063
        1013 => "0001101110",  -- +3.4578
        1014 => "0001111100",  -- +3.9032
        1015 => "0001111100",  -- +3.8784
        1016 => "0001110010",  -- +3.5815
        1017 => "0001010011",  -- +2.6166
        1018 => "0001010110",  -- +2.6908
        1019 => "0001000101",  -- +2.1713
        1020 => "0000110100",  -- +1.6270
        1021 => "0000111001",  -- +1.8002
        1022 => "0000100001",  -- +1.0579
        1023 => "0001010110",  -- +2.7156
        1024 => "0001011011",  -- +2.8640
        1025 => "0000111111",  -- +1.9981
        1026 => "0001000011",  -- +2.1218
        1027 => "0001000001",  -- +2.0476
        1028 => "0000100101",  -- +1.1816
        1029 => "0001001010",  -- +2.3197
        1030 => "0001000100",  -- +2.1465
        1031 => "0000101110",  -- +1.4538
        1032 => "0000001110",  -- +0.4394
        1033 => "0000001000",  -- +0.2662
        1034 => "1111110101",  -- -0.3276
        1035 => "0000101000",  -- +1.2806
        1036 => "0000100100",  -- +1.1321
        1037 => "0000001010",  -- +0.3157
        1038 => "0000100101",  -- +1.1569
        1039 => "0000100010",  -- +1.0827
        1040 => "1111111011",  -- -0.1297
        1041 => "0000001100",  -- +0.3899
        1042 => "0000010010",  -- +0.5631
        1043 => "1111011100",  -- -1.1193
        1044 => "0000000111",  -- +0.2415
        1045 => "0000010110",  -- +0.7115
        1046 => "1111011010",  -- -1.1688
        1047 => "0000000110",  -- +0.2167
        1048 => "0000011100",  -- +0.8847
        1049 => "1111100100",  -- -0.8472
        1050 => "0000000111",  -- +0.2415
        1051 => "0000011111",  -- +0.9837
        1052 => "1111101010",  -- -0.6740
        1053 => "0000001000",  -- +0.2662
        1054 => "0000011110",  -- +0.9590
        1055 => "1111101000",  -- -0.7482
        1056 => "0000001000",  -- +0.2662
        1057 => "0000011011",  -- +0.8600
        1058 => "1111100010",  -- -0.9214
        1059 => "0000000110",  -- +0.2167
        1060 => "0000011001",  -- +0.7858
        1061 => "1111011110",  -- -1.0451
        1062 => "0000000011",  -- +0.1177
        1063 => "0000010101",  -- +0.6868
        1064 => "1111010111",  -- -1.2678
        1065 => "1111111111",  -- -0.0307
        1066 => "0000010010",  -- +0.5631
        1067 => "1111001111",  -- -1.5152
        1068 => "1111110111",  -- -0.2534
        1069 => "0000001010",  -- +0.3404
        1070 => "1111001010",  -- -1.6636
        1071 => "1111111000",  -- -0.2286
        1072 => "0000001010",  -- +0.3157
        1073 => "1111001111",  -- -1.5152
        1074 => "0000000001",  -- +0.0435
        1075 => "0000001100",  -- +0.3899
        1076 => "1111011101",  -- -1.0698
        1077 => "1111111010",  -- -0.1791
        1078 => "1111110111",  -- -0.2534
        1079 => "1111010111",  -- -1.2678
        1080 => "0010000000",  -- +4.0269
        1081 => "0001111110",  -- +3.9526
        1082 => "0001111100",  -- +3.9032
        1083 => "0001111011",  -- +3.8537
        1084 => "0001111000",  -- +3.7547
        1085 => "0001111000",  -- +3.7547
        1086 => "0001111111",  -- +3.9774
        1087 => "0001111110",  -- +3.9526
        1088 => "0001111000",  -- +3.7547
        1089 => "0001111001",  -- +3.8042
        1090 => "0001111100",  -- +3.8784
        1091 => "0001101110",  -- +3.4578
        1092 => "0000110111",  -- +1.7259
        1093 => "0000111110",  -- +1.9486
        1094 => "0000101000",  -- +1.2558
        1095 => "0000110101",  -- +1.6764
        1096 => "0000111111",  -- +1.9733
        1097 => "0000100001",  -- +1.0332
        1098 => "0001000000",  -- +2.0228
        1099 => "0001000010",  -- +2.0723
        1100 => "0000100001",  -- +1.0332
        1101 => "0001010010",  -- +2.5919
        1102 => "0001010001",  -- +2.5424
        1103 => "0000110110",  -- +1.7012
        1104 => "0000010010",  -- +0.5631
        1105 => "0000001111",  -- +0.4889
        1106 => "1111111010",  -- -0.1791
        1107 => "0000010010",  -- +0.5878
        1108 => "0000010001",  -- +0.5384
        1109 => "1111110101",  -- -0.3276
        1110 => "0000100110",  -- +1.2064
        1111 => "0000100110",  -- +1.2064
        1112 => "1111111100",  -- -0.1049
        1113 => "0000001111",  -- +0.4889
        1114 => "0000010111",  -- +0.7363
        1115 => "1111011111",  -- -1.0203
        1116 => "0000000110",  -- +0.1920
        1117 => "0000010101",  -- +0.6868
        1118 => "1111011001",  -- -1.1935
        1119 => "0000000110",  -- +0.1920
        1120 => "0000011100",  -- +0.8847
        1121 => "1111100100",  -- -0.8719
        1122 => "0000000101",  -- +0.1672
        1123 => "0000011101",  -- +0.9342
        1124 => "1111101000",  -- -0.7482
        1125 => "0000000110",  -- +0.2167
        1126 => "0000011101",  -- +0.9342
        1127 => "1111100110",  -- -0.7977
        1128 => "0000001010",  -- +0.3157
        1129 => "0000011101",  -- +0.9342
        1130 => "1111100101",  -- -0.8224
        1131 => "0000001010",  -- +0.3404
        1132 => "0000011101",  -- +0.9095
        1133 => "1111100100",  -- -0.8719
        1134 => "0000001001",  -- +0.2909
        1135 => "0000011100",  -- +0.8847
        1136 => "1111011101",  -- -1.0698
        1137 => "0000000001",  -- +0.0435
        1138 => "0000010100",  -- +0.6373
        1139 => "1111010010",  -- -1.4162
        1140 => "1111111010",  -- -0.1791
        1141 => "0000001110",  -- +0.4394
        1142 => "1111001100",  -- -1.6141
        1143 => "1111110110",  -- -0.3029
        1144 => "0000001001",  -- +0.2909
        1145 => "1111001101",  -- -1.5894
        1146 => "1111111011",  -- -0.1297
        1147 => "0000000100",  -- +0.1425
        1148 => "1111010111",  -- -1.2678
        1149 => "1111110010",  -- -0.4266
        1150 => "1111101001",  -- -0.6987
        1151 => "1111001110",  -- -1.5399
        1152 => "0001111000",  -- +3.7795
        1153 => "0001110111",  -- +3.7300
        1154 => "0001110011",  -- +3.6063
        1155 => "0001001100",  -- +2.3939
        1156 => "0001001011",  -- +2.3692
        1157 => "0001000011",  -- +2.1218
        1158 => "0001001011",  -- +2.3692
        1159 => "0001001110",  -- +2.4682
        1160 => "0000111111",  -- +1.9981
        1161 => "0001010111",  -- +2.7403
        1162 => "0001011110",  -- +2.9630
        1163 => "0001000111",  -- +2.2455
        1164 => "0000101011",  -- +1.3548
        1165 => "0000111000",  -- +1.7507
        1166 => "0000010111",  -- +0.7363
        1167 => "0000011101",  -- +0.9342
        1168 => "0000101100",  -- +1.3796
        1169 => "0000000110",  -- +0.1920
        1170 => "0000110000",  -- +1.5033
        1171 => "0000110100",  -- +1.6270
        1172 => "0000010010",  -- +0.5878
        1173 => "0000110100",  -- +1.6270
        1174 => "0000110111",  -- +1.7259
        1175 => "0000010101",  -- +0.6868
        1176 => "0000010100",  -- +0.6373
        1177 => "0000011011",  -- +0.8600
        1178 => "1111110101",  -- -0.3276
        1179 => "0000001100",  -- +0.3899
        1180 => "0000010011",  -- +0.6126
        1181 => "1111101000",  -- -0.7482
        1182 => "0000011101",  -- +0.9342
        1183 => "0000100011",  -- +1.1074
        1184 => "1111110000",  -- -0.4760
        1185 => "0000010010",  -- +0.5878
        1186 => "0000011001",  -- +0.7858
        1187 => "1111100001",  -- -0.9461
        1188 => "0000001010",  -- +0.3404
        1189 => "0000010111",  -- +0.7363
        1190 => "1111011100",  -- -1.0946
        1191 => "0000001010",  -- +0.3157
        1192 => "0000011101",  -- +0.9095
        1193 => "1111100011",  -- -0.8966
        1194 => "0000001000",  -- +0.2662
        1195 => "0000011110",  -- +0.9590
        1196 => "1111100101",  -- -0.8224
        1197 => "0000001010",  -- +0.3157
        1198 => "0000011101",  -- +0.9342
        1199 => "1111100110",  -- -0.7977
        1200 => "0000001110",  -- +0.4394
        1201 => "0000011101",  -- +0.9095
        1202 => "1111100111",  -- -0.7729
        1203 => "0000001111",  -- +0.4889
        1204 => "0000011101",  -- +0.9095
        1205 => "1111100101",  -- -0.8224
        1206 => "0000001011",  -- +0.3652
        1207 => "0000011011",  -- +0.8600
        1208 => "1111011110",  -- -1.0451
        1209 => "0000000001",  -- +0.0435
        1210 => "0000010100",  -- +0.6373
        1211 => "1111010001",  -- -1.4409
        1212 => "1111111001",  -- -0.2039
        1213 => "0000001100",  -- +0.3899
        1214 => "1111001011",  -- -1.6389
        1215 => "1111110100",  -- -0.3523
        1216 => "0000000110",  -- +0.1920
        1217 => "1111001010",  -- -1.6636
        1218 => "1111111011",  -- -0.1544
        1219 => "1111111101",  -- -0.0802
        1220 => "1111010101",  -- -1.3172
        1221 => "1111111011",  -- -0.1297
        1222 => "1111101100",  -- -0.5997
        1223 => "1111010101",  -- -1.3172
        1224 => "0001110001",  -- +3.5320
        1225 => "0001110001",  -- +3.5568
        1226 => "0001101001",  -- +3.3094
        1227 => "0000011100",  -- +0.8847
        1228 => "0000100000",  -- +1.0084
        1229 => "0000001100",  -- +0.3899
        1230 => "0000001101",  -- +0.4146
        1231 => "0000010100",  -- +0.6373
        1232 => "1111111010",  -- -0.1791
        1233 => "0000010010",  -- +0.5878
        1234 => "0000011111",  -- +0.9837
        1235 => "1111111011",  -- -0.1297
        1236 => "0000001011",  -- +0.3652
        1237 => "0000011101",  -- +0.9095
        1238 => "1111110000",  -- -0.4760
        1239 => "0000010011",  -- +0.6126
        1240 => "0000100101",  -- +1.1816
        1241 => "1111110110",  -- -0.3029
        1242 => "0000010111",  -- +0.7363
        1243 => "0000011111",  -- +0.9837
        1244 => "1111111000",  -- -0.2286
        1245 => "0000001111",  -- +0.4889
        1246 => "0000011010",  -- +0.8352
        1247 => "1111101100",  -- -0.6245
        1248 => "0000000110",  -- +0.2167
        1249 => "0000011001",  -- +0.7858
        1250 => "1111011110",  -- -1.0451
        1251 => "0000000110",  -- +0.2167
        1252 => "0000010110",  -- +0.7115
        1253 => "1111011100",  -- -1.0946
        1254 => "0000001010",  -- +0.3404
        1255 => "0000010010",  -- +0.5878
        1256 => "1111100001",  -- -0.9461
        1257 => "0000001010",  -- +0.3157
        1258 => "0000001101",  -- +0.4146
        1259 => "1111011111",  -- -1.0203
        1260 => "0000001110",  -- +0.4641
        1261 => "0000010101",  -- +0.6868
        1262 => "1111100000",  -- -0.9709
        1263 => "0000001111",  -- +0.4889
        1264 => "0000011101",  -- +0.9342
        1265 => "1111100100",  -- -0.8719
        1266 => "0000001101",  -- +0.4146
        1267 => "0000011111",  -- +0.9837
        1268 => "1111100011",  -- -0.8966
        1269 => "0000001101",  -- +0.4146
        1270 => "0000011101",  -- +0.9095
        1271 => "1111100101",  -- -0.8224
        1272 => "0000010001",  -- +0.5384
        1273 => "0000011011",  -- +0.8600
        1274 => "1111101000",  -- -0.7235
        1275 => "0000001111",  -- +0.4889
        1276 => "0000010110",  -- +0.7115
        1277 => "1111100000",  -- -0.9709
        1278 => "0000000100",  -- +0.1425
        1279 => "0000010000",  -- +0.5136
        1280 => "1111010101",  -- -1.3420
        1281 => "1111111100",  -- -0.1049
        1282 => "0000001110",  -- +0.4394
        1283 => "1111001101",  -- -1.5647
        1284 => "1111110110",  -- -0.3029
        1285 => "0000000110",  -- +0.2167
        1286 => "1111001001",  -- -1.7131
        1287 => "1111110100",  -- -0.3523
        1288 => "1111111111",  -- -0.0060
        1289 => "1111001001",  -- -1.6884
        1290 => "1111111111",  -- -0.0060
        1291 => "1111111001",  -- -0.2039
        1292 => "1111010111",  -- -1.2678
        1293 => "0000001010",  -- +0.3404
        1294 => "1111110111",  -- -0.2534
        1295 => "1111100011",  -- -0.8966
        1296 => "0001010110",  -- +2.7156
        1297 => "0001011001",  -- +2.7898
        1298 => "0001010010",  -- +2.5671
        1299 => "0000011010",  -- +0.8352
        1300 => "0000011101",  -- +0.9342
        1301 => "0000001110",  -- +0.4641
        1302 => "0000010010",  -- +0.5878
        1303 => "0000011001",  -- +0.8105
        1304 => "0000000100",  -- +0.1425
        1305 => "0000010101",  -- +0.6868
        1306 => "0000100000",  -- +1.0084
        1307 => "0000000010",  -- +0.0930
        1308 => "0000000010",  -- +0.0683
        1309 => "0000010000",  -- +0.5136
        1310 => "1111101100",  -- -0.6245
        1311 => "1111111101",  -- -0.0802
        1312 => "0000001110",  -- +0.4394
        1313 => "1111100010",  -- -0.9214
        1314 => "1111111010",  -- -0.1791
        1315 => "0000001001",  -- +0.2909
        1316 => "1111010100",  -- -1.3667
        1317 => "1111110111",  -- -0.2781
        1318 => "0000001010",  -- +0.3157
        1319 => "1111001100",  -- -1.6141
        1320 => "1111110111",  -- -0.2534
        1321 => "0000001100",  -- +0.3899
        1322 => "1111001110",  -- -1.5399
        1323 => "1111111100",  -- -0.1049
        1324 => "0000001011",  -- +0.3652
        1325 => "1111011010",  -- -1.1688
        1326 => "1111110011",  -- -0.3771
        1327 => "1111111000",  -- -0.2286
        1328 => "1111011100",  -- -1.1193
        1329 => "1111101110",  -- -0.5503
        1330 => "1111101110",  -- -0.5503
        1331 => "1111010001",  -- -1.4409
        1332 => "0000000011",  -- +0.1177
        1333 => "0000001001",  -- +0.2909
        1334 => "1111011100",  -- -1.0946
        1335 => "0000000111",  -- +0.2415
        1336 => "0000010101",  -- +0.6621
        1337 => "1111100000",  -- -0.9709
        1338 => "0000000110",  -- +0.1920
        1339 => "0000010111",  -- +0.7363
        1340 => "1111011101",  -- -1.0698
        1341 => "0000000101",  -- +0.1672
        1342 => "0000010100",  -- +0.6373
        1343 => "1111011101",  -- -1.0698
        1344 => "0000000110",  -- +0.1920
        1345 => "0000001111",  -- +0.4889
        1346 => "1111011110",  -- -1.0451
        1347 => "0000000101",  -- +0.1672
        1348 => "0000001101",  -- +0.4146
        1349 => "1111011100",  -- -1.1193
        1350 => "0000000101",  -- +0.1672
        1351 => "0000010001",  -- +0.5384
        1352 => "1111011010",  -- -1.1688
        1353 => "0000000101",  -- +0.1672
        1354 => "0000010011",  -- +0.6126
        1355 => "1111011001",  -- -1.2183
        1356 => "0000000000",  -- +0.0188
        1357 => "0000001010",  -- +0.3404
        1358 => "1111010011",  -- -1.3915
        1359 => "1111111101",  -- -0.0802
        1360 => "1111111111",  -- -0.0307
        1361 => "1111010000",  -- -1.4904
        1362 => "0000000000",  -- +0.0188
        1363 => "1111110011",  -- -0.3771
        1364 => "1111010101",  -- -1.3420
        1365 => "0000010000",  -- +0.5136
        1366 => "1111111011",  -- -0.1544
        1367 => "1111100110",  -- -0.7977
        1368 => "0000100101",  -- +1.1816
        1369 => "0000101010",  -- +1.3301
        1370 => "0000100100",  -- +1.1321
        1371 => "0000100100",  -- +1.1321
        1372 => "0000100101",  -- +1.1569
        1373 => "0000011110",  -- +0.9590
        1374 => "0000100001",  -- +1.0579
        1375 => "0000100101",  -- +1.1569
        1376 => "0000011001",  -- +0.7858
        1377 => "0000100001",  -- +1.0332
        1378 => "0000100101",  -- +1.1816
        1379 => "0000010100",  -- +0.6373
        1380 => "0000000111",  -- +0.2415
        1381 => "0000001110",  -- +0.4641
        1382 => "1111111000",  -- -0.2286
        1383 => "1111101000",  -- -0.7235
        1384 => "1111110011",  -- -0.3771
        1385 => "1111010100",  -- -1.3667
        1386 => "1111100101",  -- -0.8224
        1387 => "1111111000",  -- -0.2286
        1388 => "1111000010",  -- -1.9110
        1389 => "1111101000",  -- -0.7482
        1390 => "1111111101",  -- -0.0802
        1391 => "1110111111",  -- -2.0100
        1392 => "1111101101",  -- -0.5750
        1393 => "1111111111",  -- -0.0060
        1394 => "1111001000",  -- -1.7378
        1395 => "1111111111",  -- -0.0307
        1396 => "0000001001",  -- +0.2909
        1397 => "1111100001",  -- -0.9461
        1398 => "0000000100",  -- +0.1425
        1399 => "0000000110",  -- +0.2167
        1400 => "1111110010",  -- -0.4266
        1401 => "1111100110",  -- -0.7977
        1402 => "1111100110",  -- -0.7977
        1403 => "1111010011",  -- -1.3915
        1404 => "1111100000",  -- -0.9709
        1405 => "1111100110",  -- -0.7977
        1406 => "1111000110",  -- -1.8121
        1407 => "1111101111",  -- -0.5255
        1408 => "1111111100",  -- -0.1049
        1409 => "1111001110",  -- -1.5399
        1410 => "1111110000",  -- -0.4760
        1411 => "0000000011",  -- +0.1177
        1412 => "1111001101",  -- -1.5894
        1413 => "1111110111",  -- -0.2534
        1414 => "0000001000",  -- +0.2662
        1415 => "1111010001",  -- -1.4409
        1416 => "0000000010",  -- +0.0930
        1417 => "0000001110",  -- +0.4641
        1418 => "1111011101",  -- -1.0698
        1419 => "0000001000",  -- +0.2662
        1420 => "0000010100",  -- +0.6373
        1421 => "1111100111",  -- -0.7729
        1422 => "0000001010",  -- +0.3404
        1423 => "0000011001",  -- +0.7858
        1424 => "1111100111",  -- -0.7729
        1425 => "0000001000",  -- +0.2662
        1426 => "0000010100",  -- +0.6373
        1427 => "1111011111",  -- -1.0203
        1428 => "0000000010",  -- +0.0683
        1429 => "0000000101",  -- +0.1672
        1430 => "1111010100",  -- -1.3667
        1431 => "1111111101",  -- -0.0802
        1432 => "1111110101",  -- -0.3276
        1433 => "1111001101",  -- -1.5894
        1434 => "0000000010",  -- +0.0930
        1435 => "1111101111",  -- -0.5008
        1436 => "1111010011",  -- -1.3915
        1437 => "0000001110",  -- +0.4641
        1438 => "1111110111",  -- -0.2534
        1439 => "1111100001",  -- -0.9461
        1440 => "0000011010",  -- +0.8352
        1441 => "0000011111",  -- +0.9837
        1442 => "0000011001",  -- +0.8105
        1443 => "0000011001",  -- +0.7858
        1444 => "0000011001",  -- +0.8105
        1445 => "0000010101",  -- +0.6868
        1446 => "0000010000",  -- +0.5136
        1447 => "0000010001",  -- +0.5384
        1448 => "0000001010",  -- +0.3404
        1449 => "0000001010",  -- +0.3157
        1450 => "0000001011",  -- +0.3652
        1451 => "0000000001",  -- +0.0435
        1452 => "0000001100",  -- +0.3899
        1453 => "0000001101",  -- +0.4146
        1454 => "1111111111",  -- -0.0060
        1455 => "1111111111",  -- -0.0060
        1456 => "0000000010",  -- +0.0930
        1457 => "1111101111",  -- -0.5008
        1458 => "1111100101",  -- -0.8224
        1459 => "1111110011",  -- -0.4018
        1460 => "1111010001",  -- -1.4657
        1461 => "1111100001",  -- -0.9461
        1462 => "1111110000",  -- -0.4760
        1463 => "1111000110",  -- -1.7873
        1464 => "1111101111",  -- -0.5255
        1465 => "1111111010",  -- -0.1791
        1466 => "1111001111",  -- -1.5152
        1467 => "0000001001",  -- +0.2909
        1468 => "0000001111",  -- +0.4889
        1469 => "1111101000",  -- -0.7235
        1470 => "0000001100",  -- +0.3899
        1471 => "0000010000",  -- +0.5136
        1472 => "1111101111",  -- -0.5255
        1473 => "1111111010",  -- -0.1791
        1474 => "1111111100",  -- -0.1049
        1475 => "1111100001",  -- -0.9461
        1476 => "1111101011",  -- -0.6492
        1477 => "1111110001",  -- -0.4513
        1478 => "1111010011",  -- -1.3915
        1479 => "1111110000",  -- -0.4760
        1480 => "1111111111",  -- -0.0060
        1481 => "1111010101",  -- -1.3420
        1482 => "1111110101",  -- -0.3276
        1483 => "0000001001",  -- +0.2909
        1484 => "1111010101",  -- -1.3420
        1485 => "1111111011",  -- -0.1297
        1486 => "0000001110",  -- +0.4394
        1487 => "1111011000",  -- -1.2430
        1488 => "0000000111",  -- +0.2415
        1489 => "0000010101",  -- +0.6868
        1490 => "1111100110",  -- -0.7977
        1491 => "0000001010",  -- +0.3157
        1492 => "0000011001",  -- +0.8105
        1493 => "1111110000",  -- -0.4760
        1494 => "0000001001",  -- +0.2909
        1495 => "0000011001",  -- +0.8105
        1496 => "1111101100",  -- -0.6245
        1497 => "0000001110",  -- +0.4641
        1498 => "0000011010",  -- +0.8352
        1499 => "1111101000",  -- -0.7235
        1500 => "0000001100",  -- +0.3899
        1501 => "0000001110",  -- +0.4394
        1502 => "1111011110",  -- -1.0451
        1503 => "1111111101",  -- -0.0802
        1504 => "1111110010",  -- -0.4266
        1505 => "1111001010",  -- -1.6636
        1506 => "0000000010",  -- +0.0683
        1507 => "1111101100",  -- -0.5997
        1508 => "1111010001",  -- -1.4657
        1509 => "0000000110",  -- +0.2167
        1510 => "1111101110",  -- -0.5503
        1511 => "1111011000",  -- -1.2430
        1512 => "0000001000",  -- +0.2662
        1513 => "0000001100",  -- +0.3899
        1514 => "0000000011",  -- +0.1177
        1515 => "0000000101",  -- +0.1672
        1516 => "0000000101",  -- +0.1672
        1517 => "1111111110",  -- -0.0554
        1518 => "0000001001",  -- +0.2909
        1519 => "0000001000",  -- +0.2662
        1520 => "0000000000",  -- +0.0188
        1521 => "0000001110",  -- +0.4641
        1522 => "0000001100",  -- +0.3899
        1523 => "0000000010",  -- +0.0683
        1524 => "0000010101",  -- +0.6621
        1525 => "0000010001",  -- +0.5384
        1526 => "0000000100",  -- +0.1425
        1527 => "0000010111",  -- +0.7363
        1528 => "0000010011",  -- +0.6126
        1529 => "0000000110",  -- +0.1920
        1530 => "0000001010",  -- +0.3157
        1531 => "0000001100",  -- +0.3899
        1532 => "1111111100",  -- -0.1049
        1533 => "1111111011",  -- -0.1297
        1534 => "1111111101",  -- -0.0802
        1535 => "1111101001",  -- -0.6987
        1536 => "0000000010",  -- +0.0683
        1537 => "0000000001",  -- +0.0435
        1538 => "1111100100",  -- -0.8472
        1539 => "0000001000",  -- +0.2662
        1540 => "0000001010",  -- +0.3404
        1541 => "1111100100",  -- -0.8472
        1542 => "0000000011",  -- +0.1177
        1543 => "0000001010",  -- +0.3404
        1544 => "1111011101",  -- -1.0698
        1545 => "1111111111",  -- -0.0307
        1546 => "0000000101",  -- +0.1672
        1547 => "1111011111",  -- -1.0203
        1548 => "1111110011",  -- -0.4018
        1549 => "1111111011",  -- -0.1544
        1550 => "1111011000",  -- -1.2430
        1551 => "1111110011",  -- -0.3771
        1552 => "0000000011",  -- +0.1177
        1553 => "1111010101",  -- -1.3172
        1554 => "1111111001",  -- -0.2039
        1555 => "0000001110",  -- +0.4394
        1556 => "1111011001",  -- -1.1935
        1557 => "1111111111",  -- -0.0060
        1558 => "0000010010",  -- +0.5878
        1559 => "1111011110",  -- -1.0451
        1560 => "0000010010",  -- +0.5878
        1561 => "0000100010",  -- +1.0827
        1562 => "1111110100",  -- -0.3523
        1563 => "0000010110",  -- +0.7115
        1564 => "0000101000",  -- +1.2806
        1565 => "0000000000",  -- +0.0188
        1566 => "0000001011",  -- +0.3652
        1567 => "0000011111",  -- +0.9837
        1568 => "1111110001",  -- -0.4513
        1569 => "0000001001",  -- +0.2909
        1570 => "0000011001",  -- +0.7858
        1571 => "1111100101",  -- -0.8224
        1572 => "0000010000",  -- +0.5136
        1573 => "0000010110",  -- +0.7115
        1574 => "1111100011",  -- -0.8966
        1575 => "0000001101",  -- +0.4146
        1576 => "0000000111",  -- +0.2415
        1577 => "1111011011",  -- -1.1441
        1578 => "0000000010",  -- +0.0930
        1579 => "1111101111",  -- -0.5255
        1580 => "1111001111",  -- -1.5152
        1581 => "0000000110",  -- +0.1920
        1582 => "1111101011",  -- -0.6492
        1583 => "1111010100",  -- -1.3667
        1584 => "0000000110",  -- +0.2167
        1585 => "0000001000",  -- +0.2662
        1586 => "1111111100",  -- -0.1049
        1587 => "0000001100",  -- +0.3899
        1588 => "0000001101",  -- +0.4146
        1589 => "1111111110",  -- -0.0554
        1590 => "0000010000",  -- +0.5136
        1591 => "0000001111",  -- +0.4889
        1592 => "0000000000",  -- +0.0188
        1593 => "0000010010",  -- +0.5631
        1594 => "0000001101",  -- +0.4146
        1595 => "1111111110",  -- -0.0554
        1596 => "0000010001",  -- +0.5384
        1597 => "0000001010",  -- +0.3157
        1598 => "1111111010",  -- -0.1791
        1599 => "0000001010",  -- +0.3404
        1600 => "0000000010",  -- +0.0683
        1601 => "1111110010",  -- -0.4266
        1602 => "0000000101",  -- +0.1672
        1603 => "1111111100",  -- -0.1049
        1604 => "1111101110",  -- -0.5503
        1605 => "0000000011",  -- +0.1177
        1606 => "1111111000",  -- -0.2286
        1607 => "1111101001",  -- -0.6987
        1608 => "1111110111",  -- -0.2534
        1609 => "1111101100",  -- -0.5997
        1610 => "1111011000",  -- -1.2430
        1611 => "1111110100",  -- -0.3523
        1612 => "1111110001",  -- -0.4513
        1613 => "1111010100",  -- -1.3667
        1614 => "1111111011",  -- -0.1544
        1615 => "0000000010",  -- +0.0683
        1616 => "1111011011",  -- -1.1441
        1617 => "0000000001",  -- +0.0435
        1618 => "0000001010",  -- +0.3404
        1619 => "1111100001",  -- -0.9461
        1620 => "1111111000",  -- -0.2286
        1621 => "0000000010",  -- +0.0930
        1622 => "1111011000",  -- -1.2430
        1623 => "1111110001",  -- -0.4513
        1624 => "0000000011",  -- +0.1177
        1625 => "1111010000",  -- -1.4904
        1626 => "1111110111",  -- -0.2781
        1627 => "0000001101",  -- +0.4146
        1628 => "1111010111",  -- -1.2678
        1629 => "1111111111",  -- -0.0307
        1630 => "0000010010",  -- +0.5631
        1631 => "1111011111",  -- -1.0203
        1632 => "0000010101",  -- +0.6621
        1633 => "0000100101",  -- +1.1569
        1634 => "1111111000",  -- -0.2286
        1635 => "0000011001",  -- +0.8105
        1636 => "0000101101",  -- +1.4290
        1637 => "0000000011",  -- +0.1177
        1638 => "0000001011",  -- +0.3652
        1639 => "0000100001",  -- +1.0579
        1640 => "1111110000",  -- -0.4760
        1641 => "0000000010",  -- +0.0930
        1642 => "0000011001",  -- +0.7858
        1643 => "1111100000",  -- -0.9956
        1644 => "0000000100",  -- +0.1425
        1645 => "0000010010",  -- +0.5878
        1646 => "1111011001",  -- -1.2183
        1647 => "0000001010",  -- +0.3157
        1648 => "0000001101",  -- +0.4146
        1649 => "1111011001",  -- -1.1935
        1650 => "0000001010",  -- +0.3157
        1651 => "1111111000",  -- -0.2286
        1652 => "1111010101",  -- -1.3172
        1653 => "0000001000",  -- +0.2662
        1654 => "1111101100",  -- -0.5997
        1655 => "1111010100",  -- -1.3667
        1656 => "0000001110",  -- +0.4394
        1657 => "0000001101",  -- +0.4146
        1658 => "1111111101",  -- -0.0802
        1659 => "0000001111",  -- +0.4889
        1660 => "0000001110",  -- +0.4394
        1661 => "1111111010",  -- -0.1791
        1662 => "0000001101",  -- +0.4146
        1663 => "0000001000",  -- +0.2662
        1664 => "1111110100",  -- -0.3523
        1665 => "0000000111",  -- +0.2415
        1666 => "1111111101",  -- -0.0802
        1667 => "1111101011",  -- -0.6492
        1668 => "0000000000",  -- +0.0188
        1669 => "1111110010",  -- -0.4266
        1670 => "1111100000",  -- -0.9709
        1671 => "1111111000",  -- -0.2286
        1672 => "1111101000",  -- -0.7482
        1673 => "1111010111",  -- -1.2678
        1674 => "1111111100",  -- -0.1049
        1675 => "1111101100",  -- -0.6245
        1676 => "1111011001",  -- -1.1935
        1677 => "0000001010",  -- +0.3404
        1678 => "1111111010",  -- -0.1791
        1679 => "1111100111",  -- -0.7729
        1680 => "0000000010",  -- +0.0683
        1681 => "1111110011",  -- -0.4018
        1682 => "1111100000",  -- -0.9956
        1683 => "1111110010",  -- -0.4266
        1684 => "1111101010",  -- -0.6740
        1685 => "1111010011",  -- -1.3915
        1686 => "1111110100",  -- -0.3523
        1687 => "1111110110",  -- -0.3029
        1688 => "1111011001",  -- -1.2183
        1689 => "0000000001",  -- +0.0435
        1690 => "0000000010",  -- +0.0930
        1691 => "1111011111",  -- -1.0203
        1692 => "1111111110",  -- -0.0554
        1693 => "1111111111",  -- -0.0307
        1694 => "1111010110",  -- -1.2925
        1695 => "1111110101",  -- -0.3276
        1696 => "1111111101",  -- -0.0802
        1697 => "1111010000",  -- -1.4904
        1698 => "1111110111",  -- -0.2781
        1699 => "0000000011",  -- +0.1177
        1700 => "1111010101",  -- -1.3420
        1701 => "1111110111",  -- -0.2781
        1702 => "0000000010",  -- +0.0683
        1703 => "1111010111",  -- -1.2678
        1704 => "0000000000",  -- +0.0188
        1705 => "0000001011",  -- +0.3652
        1706 => "1111100100",  -- -0.8719
        1707 => "0000000111",  -- +0.2415
        1708 => "0000011001",  -- +0.8105
        1709 => "1111101111",  -- -0.5255
        1710 => "0000000010",  -- +0.0683
        1711 => "0000011001",  -- +0.7858
        1712 => "1111101000",  -- -0.7482
        1713 => "1111111100",  -- -0.1049
        1714 => "0000010010",  -- +0.5878
        1715 => "1111011100",  -- -1.1193
        1716 => "1111111101",  -- -0.0802
        1717 => "0000001110",  -- +0.4641
        1718 => "1111010110",  -- -1.2925
        1719 => "0000000001",  -- +0.0435
        1720 => "0000001010",  -- +0.3404
        1721 => "1111010110",  -- -1.2925
        1722 => "0000000101",  -- +0.1672
        1723 => "1111110110",  -- -0.3029
        1724 => "1111010011",  -- -1.3915
        1725 => "0000000100",  -- +0.1425
        1726 => "1111100111",  -- -0.7729
        1727 => "1111001111"   -- -1.5152
    );
    
begin
    
    process(clk)
    begin
        if rising_edge(clk) then
            if re = '1' then
                dout_reg <= mem(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

    -- Output assignment
    dout <= dout_reg;
end architecture rtl;
