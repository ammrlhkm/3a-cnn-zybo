--------------------------------------------------------------------------------
-- VHDL ROM with grayscale image pixel initialization (Read-Only)
-- Generated from: tiger_320x240.ppm
-- Generated on: 2025-12-18 17:14:14
-- Image size: 320x240 Grayscale
-- Memory depth: 76800 bytes
-- Address bits: 17
-- Conversion: Y = 0.299*R + 0.587*G + 0.114*B
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity disp_input_rom is
    generic (
        CELL_COUNT : integer := 76800;
        ADDR_WIDTH : integer := 17;
        DATA_WIDTH : integer := 8
    );
    port (
        clk     : in  std_logic;
        addr    : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        re      : in  std_logic;
        dout    : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end entity disp_input_rom;

architecture rtl of disp_input_rom is
    
    -- Memory type
    type mem_type is array (0 to 76799) of std_logic_vector(DATA_WIDTH-1 downto 0);

    -- Output register for better timing (addresses SYNTH-6 warning)
    signal dout_reg : std_logic_vector(DATA_WIDTH-1 downto 0) := (others => '0');

    -- Constant memory with grayscale pixels
    constant mem : mem_type := (
        0 => X"3E",  -- 62
        1 => X"3E",  -- 62
        2 => X"3D",  -- 61
        3 => X"3D",  -- 61
        4 => X"3C",  -- 60
        5 => X"3D",  -- 61
        6 => X"3E",  -- 62
        7 => X"3E",  -- 62
        8 => X"3D",  -- 61
        9 => X"3D",  -- 61
        10 => X"3D",  -- 61
        11 => X"3E",  -- 62
        12 => X"3F",  -- 63
        13 => X"41",  -- 65
        14 => X"43",  -- 67
        15 => X"44",  -- 68
        16 => X"43",  -- 67
        17 => X"43",  -- 67
        18 => X"43",  -- 67
        19 => X"44",  -- 68
        20 => X"44",  -- 68
        21 => X"44",  -- 68
        22 => X"44",  -- 68
        23 => X"45",  -- 69
        24 => X"46",  -- 70
        25 => X"47",  -- 71
        26 => X"47",  -- 71
        27 => X"47",  -- 71
        28 => X"47",  -- 71
        29 => X"46",  -- 70
        30 => X"45",  -- 69
        31 => X"45",  -- 69
        32 => X"44",  -- 68
        33 => X"44",  -- 68
        34 => X"43",  -- 67
        35 => X"42",  -- 66
        36 => X"42",  -- 66
        37 => X"42",  -- 66
        38 => X"41",  -- 65
        39 => X"41",  -- 65
        40 => X"40",  -- 64
        41 => X"3F",  -- 63
        42 => X"3D",  -- 61
        43 => X"3C",  -- 60
        44 => X"3B",  -- 59
        45 => X"3A",  -- 58
        46 => X"39",  -- 57
        47 => X"39",  -- 57
        48 => X"38",  -- 56
        49 => X"38",  -- 56
        50 => X"37",  -- 55
        51 => X"36",  -- 54
        52 => X"35",  -- 53
        53 => X"35",  -- 53
        54 => X"34",  -- 52
        55 => X"34",  -- 52
        56 => X"34",  -- 52
        57 => X"33",  -- 51
        58 => X"32",  -- 50
        59 => X"32",  -- 50
        60 => X"32",  -- 50
        61 => X"33",  -- 51
        62 => X"34",  -- 52
        63 => X"35",  -- 53
        64 => X"36",  -- 54
        65 => X"38",  -- 56
        66 => X"3A",  -- 58
        67 => X"3C",  -- 60
        68 => X"3D",  -- 61
        69 => X"3F",  -- 63
        70 => X"43",  -- 67
        71 => X"45",  -- 69
        72 => X"48",  -- 72
        73 => X"49",  -- 73
        74 => X"4B",  -- 75
        75 => X"4D",  -- 77
        76 => X"4E",  -- 78
        77 => X"4F",  -- 79
        78 => X"4E",  -- 78
        79 => X"4E",  -- 78
        80 => X"4F",  -- 79
        81 => X"4E",  -- 78
        82 => X"4E",  -- 78
        83 => X"4F",  -- 79
        84 => X"4E",  -- 78
        85 => X"4F",  -- 79
        86 => X"4E",  -- 78
        87 => X"4E",  -- 78
        88 => X"51",  -- 81
        89 => X"4C",  -- 76
        90 => X"4C",  -- 76
        91 => X"54",  -- 84
        92 => X"66",  -- 102
        93 => X"7A",  -- 122
        94 => X"86",  -- 134
        95 => X"8D",  -- 141
        96 => X"8F",  -- 143
        97 => X"95",  -- 149
        98 => X"96",  -- 150
        99 => X"8D",  -- 141
        100 => X"8B",  -- 139
        101 => X"8D",  -- 141
        102 => X"8C",  -- 140
        103 => X"84",  -- 132
        104 => X"82",  -- 130
        105 => X"63",  -- 99
        106 => X"52",  -- 82
        107 => X"4E",  -- 78
        108 => X"47",  -- 71
        109 => X"48",  -- 72
        110 => X"47",  -- 71
        111 => X"38",  -- 56
        112 => X"3D",  -- 61
        113 => X"56",  -- 86
        114 => X"75",  -- 117
        115 => X"83",  -- 131
        116 => X"89",  -- 137
        117 => X"96",  -- 150
        118 => X"95",  -- 149
        119 => X"82",  -- 130
        120 => X"85",  -- 133
        121 => X"70",  -- 112
        122 => X"5A",  -- 90
        123 => X"54",  -- 84
        124 => X"52",  -- 82
        125 => X"45",  -- 69
        126 => X"42",  -- 66
        127 => X"4E",  -- 78
        128 => X"41",  -- 65
        129 => X"58",  -- 88
        130 => X"66",  -- 102
        131 => X"74",  -- 116
        132 => X"7A",  -- 122
        133 => X"80",  -- 128
        134 => X"98",  -- 152
        135 => X"A2",  -- 162
        136 => X"AA",  -- 170
        137 => X"A8",  -- 168
        138 => X"A9",  -- 169
        139 => X"AC",  -- 172
        140 => X"AE",  -- 174
        141 => X"B0",  -- 176
        142 => X"B0",  -- 176
        143 => X"AF",  -- 175
        144 => X"AE",  -- 174
        145 => X"A3",  -- 163
        146 => X"A8",  -- 168
        147 => X"AC",  -- 172
        148 => X"A5",  -- 165
        149 => X"A7",  -- 167
        150 => X"AA",  -- 170
        151 => X"9F",  -- 159
        152 => X"A0",  -- 160
        153 => X"9F",  -- 159
        154 => X"A2",  -- 162
        155 => X"9A",  -- 154
        156 => X"85",  -- 133
        157 => X"71",  -- 113
        158 => X"60",  -- 96
        159 => X"4A",  -- 74
        160 => X"45",  -- 69
        161 => X"3D",  -- 61
        162 => X"3A",  -- 58
        163 => X"3D",  -- 61
        164 => X"43",  -- 67
        165 => X"4D",  -- 77
        166 => X"5F",  -- 95
        167 => X"72",  -- 114
        168 => X"75",  -- 117
        169 => X"76",  -- 118
        170 => X"77",  -- 119
        171 => X"78",  -- 120
        172 => X"79",  -- 121
        173 => X"7B",  -- 123
        174 => X"7D",  -- 125
        175 => X"7F",  -- 127
        176 => X"7F",  -- 127
        177 => X"82",  -- 130
        178 => X"88",  -- 136
        179 => X"8C",  -- 140
        180 => X"8D",  -- 141
        181 => X"8C",  -- 140
        182 => X"8D",  -- 141
        183 => X"8C",  -- 140
        184 => X"8F",  -- 143
        185 => X"8B",  -- 139
        186 => X"87",  -- 135
        187 => X"80",  -- 128
        188 => X"71",  -- 113
        189 => X"68",  -- 104
        190 => X"70",  -- 112
        191 => X"81",  -- 129
        192 => X"8D",  -- 141
        193 => X"94",  -- 148
        194 => X"9E",  -- 158
        195 => X"A4",  -- 164
        196 => X"A5",  -- 165
        197 => X"A7",  -- 167
        198 => X"AC",  -- 172
        199 => X"B0",  -- 176
        200 => X"B0",  -- 176
        201 => X"B2",  -- 178
        202 => X"B4",  -- 180
        203 => X"B2",  -- 178
        204 => X"AE",  -- 174
        205 => X"AC",  -- 172
        206 => X"AD",  -- 173
        207 => X"AF",  -- 175
        208 => X"B5",  -- 181
        209 => X"B3",  -- 179
        210 => X"B2",  -- 178
        211 => X"B5",  -- 181
        212 => X"B8",  -- 184
        213 => X"BA",  -- 186
        214 => X"B7",  -- 183
        215 => X"B3",  -- 179
        216 => X"AF",  -- 175
        217 => X"B3",  -- 179
        218 => X"B5",  -- 181
        219 => X"B0",  -- 176
        220 => X"A9",  -- 169
        221 => X"A4",  -- 164
        222 => X"A5",  -- 165
        223 => X"A6",  -- 166
        224 => X"A6",  -- 166
        225 => X"A1",  -- 161
        226 => X"9E",  -- 158
        227 => X"A0",  -- 160
        228 => X"A2",  -- 162
        229 => X"A1",  -- 161
        230 => X"A2",  -- 162
        231 => X"A6",  -- 166
        232 => X"A3",  -- 163
        233 => X"A1",  -- 161
        234 => X"A0",  -- 160
        235 => X"A0",  -- 160
        236 => X"A2",  -- 162
        237 => X"A4",  -- 164
        238 => X"A4",  -- 164
        239 => X"A3",  -- 163
        240 => X"AB",  -- 171
        241 => X"AC",  -- 172
        242 => X"AF",  -- 175
        243 => X"B0",  -- 176
        244 => X"AF",  -- 175
        245 => X"B0",  -- 176
        246 => X"B2",  -- 178
        247 => X"B4",  -- 180
        248 => X"B0",  -- 176
        249 => X"B2",  -- 178
        250 => X"B4",  -- 180
        251 => X"AF",  -- 175
        252 => X"A5",  -- 165
        253 => X"9B",  -- 155
        254 => X"93",  -- 147
        255 => X"90",  -- 144
        256 => X"8B",  -- 139
        257 => X"92",  -- 146
        258 => X"94",  -- 148
        259 => X"8D",  -- 141
        260 => X"7D",  -- 125
        261 => X"6E",  -- 110
        262 => X"69",  -- 105
        263 => X"68",  -- 104
        264 => X"54",  -- 84
        265 => X"58",  -- 88
        266 => X"5E",  -- 94
        267 => X"5C",  -- 92
        268 => X"57",  -- 87
        269 => X"58",  -- 88
        270 => X"65",  -- 101
        271 => X"73",  -- 115
        272 => X"83",  -- 131
        273 => X"95",  -- 149
        274 => X"9E",  -- 158
        275 => X"9F",  -- 159
        276 => X"A6",  -- 166
        277 => X"A8",  -- 168
        278 => X"AA",  -- 170
        279 => X"B1",  -- 177
        280 => X"B8",  -- 184
        281 => X"B8",  -- 184
        282 => X"B7",  -- 183
        283 => X"B5",  -- 181
        284 => X"B4",  -- 180
        285 => X"B5",  -- 181
        286 => X"B8",  -- 184
        287 => X"BB",  -- 187
        288 => X"B9",  -- 185
        289 => X"BD",  -- 189
        290 => X"C1",  -- 193
        291 => X"C0",  -- 192
        292 => X"BC",  -- 188
        293 => X"BA",  -- 186
        294 => X"BD",  -- 189
        295 => X"C0",  -- 192
        296 => X"BD",  -- 189
        297 => X"BF",  -- 191
        298 => X"C0",  -- 192
        299 => X"BF",  -- 191
        300 => X"BC",  -- 188
        301 => X"BA",  -- 186
        302 => X"BA",  -- 186
        303 => X"BB",  -- 187
        304 => X"BA",  -- 186
        305 => X"B8",  -- 184
        306 => X"B6",  -- 182
        307 => X"B7",  -- 183
        308 => X"BA",  -- 186
        309 => X"BD",  -- 189
        310 => X"BF",  -- 191
        311 => X"C0",  -- 192
        312 => X"BC",  -- 188
        313 => X"BC",  -- 188
        314 => X"BE",  -- 190
        315 => X"BF",  -- 191
        316 => X"BE",  -- 190
        317 => X"BA",  -- 186
        318 => X"B2",  -- 178
        319 => X"AD",  -- 173
        320 => X"33",  -- 51
        321 => X"33",  -- 51
        322 => X"32",  -- 50
        323 => X"32",  -- 50
        324 => X"31",  -- 49
        325 => X"32",  -- 50
        326 => X"32",  -- 50
        327 => X"33",  -- 51
        328 => X"32",  -- 50
        329 => X"32",  -- 50
        330 => X"32",  -- 50
        331 => X"33",  -- 51
        332 => X"34",  -- 52
        333 => X"36",  -- 54
        334 => X"38",  -- 56
        335 => X"39",  -- 57
        336 => X"39",  -- 57
        337 => X"39",  -- 57
        338 => X"39",  -- 57
        339 => X"39",  -- 57
        340 => X"3A",  -- 58
        341 => X"3A",  -- 58
        342 => X"3A",  -- 58
        343 => X"3A",  -- 58
        344 => X"3B",  -- 59
        345 => X"3B",  -- 59
        346 => X"3C",  -- 60
        347 => X"3C",  -- 60
        348 => X"3B",  -- 59
        349 => X"3B",  -- 59
        350 => X"3A",  -- 58
        351 => X"39",  -- 57
        352 => X"38",  -- 56
        353 => X"38",  -- 56
        354 => X"38",  -- 56
        355 => X"37",  -- 55
        356 => X"37",  -- 55
        357 => X"36",  -- 54
        358 => X"36",  -- 54
        359 => X"35",  -- 53
        360 => X"34",  -- 52
        361 => X"34",  -- 52
        362 => X"32",  -- 50
        363 => X"31",  -- 49
        364 => X"30",  -- 48
        365 => X"2F",  -- 47
        366 => X"2E",  -- 46
        367 => X"2E",  -- 46
        368 => X"2C",  -- 44
        369 => X"2C",  -- 44
        370 => X"2C",  -- 44
        371 => X"2B",  -- 43
        372 => X"2A",  -- 42
        373 => X"29",  -- 41
        374 => X"29",  -- 41
        375 => X"28",  -- 40
        376 => X"28",  -- 40
        377 => X"27",  -- 39
        378 => X"26",  -- 38
        379 => X"26",  -- 38
        380 => X"26",  -- 38
        381 => X"27",  -- 39
        382 => X"28",  -- 40
        383 => X"29",  -- 41
        384 => X"2A",  -- 42
        385 => X"2C",  -- 44
        386 => X"2F",  -- 47
        387 => X"30",  -- 48
        388 => X"32",  -- 50
        389 => X"34",  -- 52
        390 => X"37",  -- 55
        391 => X"39",  -- 57
        392 => X"3C",  -- 60
        393 => X"3E",  -- 62
        394 => X"40",  -- 64
        395 => X"41",  -- 65
        396 => X"43",  -- 67
        397 => X"43",  -- 67
        398 => X"43",  -- 67
        399 => X"43",  -- 67
        400 => X"43",  -- 67
        401 => X"43",  -- 67
        402 => X"43",  -- 67
        403 => X"44",  -- 68
        404 => X"43",  -- 67
        405 => X"44",  -- 68
        406 => X"43",  -- 67
        407 => X"44",  -- 68
        408 => X"47",  -- 71
        409 => X"45",  -- 69
        410 => X"47",  -- 71
        411 => X"50",  -- 80
        412 => X"61",  -- 97
        413 => X"72",  -- 114
        414 => X"7E",  -- 126
        415 => X"83",  -- 131
        416 => X"84",  -- 132
        417 => X"88",  -- 136
        418 => X"88",  -- 136
        419 => X"84",  -- 132
        420 => X"83",  -- 131
        421 => X"86",  -- 134
        422 => X"81",  -- 129
        423 => X"78",  -- 120
        424 => X"74",  -- 116
        425 => X"56",  -- 86
        426 => X"48",  -- 72
        427 => X"4C",  -- 76
        428 => X"4C",  -- 76
        429 => X"41",  -- 65
        430 => X"34",  -- 52
        431 => X"2A",  -- 42
        432 => X"34",  -- 52
        433 => X"50",  -- 80
        434 => X"6B",  -- 107
        435 => X"74",  -- 116
        436 => X"7B",  -- 123
        437 => X"83",  -- 131
        438 => X"7D",  -- 125
        439 => X"73",  -- 115
        440 => X"7F",  -- 127
        441 => X"6B",  -- 107
        442 => X"59",  -- 89
        443 => X"4C",  -- 76
        444 => X"42",  -- 66
        445 => X"39",  -- 57
        446 => X"3B",  -- 59
        447 => X"3F",  -- 63
        448 => X"38",  -- 56
        449 => X"57",  -- 87
        450 => X"6B",  -- 107
        451 => X"7C",  -- 124
        452 => X"80",  -- 128
        453 => X"84",  -- 132
        454 => X"9C",  -- 156
        455 => X"A5",  -- 165
        456 => X"A6",  -- 166
        457 => X"A4",  -- 164
        458 => X"A6",  -- 166
        459 => X"A7",  -- 167
        460 => X"A9",  -- 169
        461 => X"A9",  -- 169
        462 => X"A8",  -- 168
        463 => X"A6",  -- 166
        464 => X"A3",  -- 163
        465 => X"9C",  -- 156
        466 => X"A3",  -- 163
        467 => X"A9",  -- 169
        468 => X"A1",  -- 161
        469 => X"A3",  -- 163
        470 => X"A5",  -- 165
        471 => X"9B",  -- 155
        472 => X"9E",  -- 158
        473 => X"A1",  -- 161
        474 => X"A5",  -- 165
        475 => X"94",  -- 148
        476 => X"76",  -- 118
        477 => X"62",  -- 98
        478 => X"58",  -- 88
        479 => X"4F",  -- 79
        480 => X"3F",  -- 63
        481 => X"41",  -- 65
        482 => X"3E",  -- 62
        483 => X"3B",  -- 59
        484 => X"3D",  -- 61
        485 => X"4B",  -- 75
        486 => X"5E",  -- 94
        487 => X"6B",  -- 107
        488 => X"72",  -- 114
        489 => X"73",  -- 115
        490 => X"76",  -- 118
        491 => X"78",  -- 120
        492 => X"7A",  -- 122
        493 => X"7E",  -- 126
        494 => X"83",  -- 131
        495 => X"85",  -- 133
        496 => X"84",  -- 132
        497 => X"85",  -- 133
        498 => X"88",  -- 136
        499 => X"89",  -- 137
        500 => X"89",  -- 137
        501 => X"89",  -- 137
        502 => X"8A",  -- 138
        503 => X"8C",  -- 140
        504 => X"8B",  -- 139
        505 => X"8C",  -- 140
        506 => X"8D",  -- 141
        507 => X"8E",  -- 142
        508 => X"83",  -- 131
        509 => X"78",  -- 120
        510 => X"7B",  -- 123
        511 => X"86",  -- 134
        512 => X"93",  -- 147
        513 => X"99",  -- 153
        514 => X"A0",  -- 160
        515 => X"A4",  -- 164
        516 => X"A4",  -- 164
        517 => X"A6",  -- 166
        518 => X"AA",  -- 170
        519 => X"AF",  -- 175
        520 => X"AF",  -- 175
        521 => X"B0",  -- 176
        522 => X"B0",  -- 176
        523 => X"AE",  -- 174
        524 => X"AB",  -- 171
        525 => X"AA",  -- 170
        526 => X"AB",  -- 171
        527 => X"AB",  -- 171
        528 => X"AE",  -- 174
        529 => X"AC",  -- 172
        530 => X"AA",  -- 170
        531 => X"AC",  -- 172
        532 => X"B0",  -- 176
        533 => X"B3",  -- 179
        534 => X"B1",  -- 177
        535 => X"AF",  -- 175
        536 => X"A8",  -- 168
        537 => X"AA",  -- 170
        538 => X"AD",  -- 173
        539 => X"AA",  -- 170
        540 => X"A6",  -- 166
        541 => X"A3",  -- 163
        542 => X"A3",  -- 163
        543 => X"A3",  -- 163
        544 => X"9A",  -- 154
        545 => X"98",  -- 152
        546 => X"98",  -- 152
        547 => X"9D",  -- 157
        548 => X"9E",  -- 158
        549 => X"9B",  -- 155
        550 => X"97",  -- 151
        551 => X"98",  -- 152
        552 => X"9F",  -- 159
        553 => X"9E",  -- 158
        554 => X"9D",  -- 157
        555 => X"9E",  -- 158
        556 => X"9F",  -- 159
        557 => X"A0",  -- 160
        558 => X"A0",  -- 160
        559 => X"9E",  -- 158
        560 => X"A2",  -- 162
        561 => X"A4",  -- 164
        562 => X"A7",  -- 167
        563 => X"A8",  -- 168
        564 => X"A8",  -- 168
        565 => X"A9",  -- 169
        566 => X"AC",  -- 172
        567 => X"AE",  -- 174
        568 => X"AC",  -- 172
        569 => X"AE",  -- 174
        570 => X"B0",  -- 176
        571 => X"AE",  -- 174
        572 => X"A6",  -- 166
        573 => X"9C",  -- 156
        574 => X"92",  -- 146
        575 => X"8C",  -- 140
        576 => X"89",  -- 137
        577 => X"8D",  -- 141
        578 => X"90",  -- 144
        579 => X"89",  -- 137
        580 => X"7D",  -- 125
        581 => X"6E",  -- 110
        582 => X"65",  -- 101
        583 => X"5F",  -- 95
        584 => X"50",  -- 80
        585 => X"52",  -- 82
        586 => X"51",  -- 81
        587 => X"4C",  -- 76
        588 => X"4C",  -- 76
        589 => X"53",  -- 83
        590 => X"5E",  -- 94
        591 => X"66",  -- 102
        592 => X"6F",  -- 111
        593 => X"81",  -- 129
        594 => X"8A",  -- 138
        595 => X"92",  -- 146
        596 => X"A0",  -- 160
        597 => X"A7",  -- 167
        598 => X"A7",  -- 167
        599 => X"AD",  -- 173
        600 => X"AE",  -- 174
        601 => X"B1",  -- 177
        602 => X"B3",  -- 179
        603 => X"B5",  -- 181
        604 => X"B4",  -- 180
        605 => X"B3",  -- 179
        606 => X"B3",  -- 179
        607 => X"B4",  -- 180
        608 => X"B8",  -- 184
        609 => X"B9",  -- 185
        610 => X"BA",  -- 186
        611 => X"BB",  -- 187
        612 => X"BC",  -- 188
        613 => X"BB",  -- 187
        614 => X"BA",  -- 186
        615 => X"B9",  -- 185
        616 => X"BC",  -- 188
        617 => X"BC",  -- 188
        618 => X"BB",  -- 187
        619 => X"BA",  -- 186
        620 => X"B8",  -- 184
        621 => X"B6",  -- 182
        622 => X"B5",  -- 181
        623 => X"B4",  -- 180
        624 => X"B7",  -- 183
        625 => X"B6",  -- 182
        626 => X"B5",  -- 181
        627 => X"B6",  -- 182
        628 => X"B7",  -- 183
        629 => X"B8",  -- 184
        630 => X"B6",  -- 182
        631 => X"B5",  -- 181
        632 => X"B8",  -- 184
        633 => X"B8",  -- 184
        634 => X"BA",  -- 186
        635 => X"BC",  -- 188
        636 => X"BC",  -- 188
        637 => X"B8",  -- 184
        638 => X"B1",  -- 177
        639 => X"AC",  -- 172
        640 => X"31",  -- 49
        641 => X"31",  -- 49
        642 => X"30",  -- 48
        643 => X"30",  -- 48
        644 => X"2F",  -- 47
        645 => X"2F",  -- 47
        646 => X"30",  -- 48
        647 => X"30",  -- 48
        648 => X"2F",  -- 47
        649 => X"2F",  -- 47
        650 => X"2F",  -- 47
        651 => X"30",  -- 48
        652 => X"31",  -- 49
        653 => X"33",  -- 51
        654 => X"35",  -- 53
        655 => X"36",  -- 54
        656 => X"37",  -- 55
        657 => X"37",  -- 55
        658 => X"37",  -- 55
        659 => X"37",  -- 55
        660 => X"37",  -- 55
        661 => X"38",  -- 56
        662 => X"38",  -- 56
        663 => X"38",  -- 56
        664 => X"38",  -- 56
        665 => X"38",  -- 56
        666 => X"38",  -- 56
        667 => X"38",  -- 56
        668 => X"38",  -- 56
        669 => X"37",  -- 55
        670 => X"37",  -- 55
        671 => X"36",  -- 54
        672 => X"35",  -- 53
        673 => X"35",  -- 53
        674 => X"34",  -- 52
        675 => X"33",  -- 51
        676 => X"34",  -- 52
        677 => X"33",  -- 51
        678 => X"32",  -- 50
        679 => X"32",  -- 50
        680 => X"31",  -- 49
        681 => X"30",  -- 48
        682 => X"2F",  -- 47
        683 => X"2E",  -- 46
        684 => X"2C",  -- 44
        685 => X"2B",  -- 43
        686 => X"2B",  -- 43
        687 => X"2A",  -- 42
        688 => X"29",  -- 41
        689 => X"29",  -- 41
        690 => X"28",  -- 40
        691 => X"27",  -- 39
        692 => X"27",  -- 39
        693 => X"26",  -- 38
        694 => X"25",  -- 37
        695 => X"25",  -- 37
        696 => X"23",  -- 35
        697 => X"22",  -- 34
        698 => X"21",  -- 33
        699 => X"21",  -- 33
        700 => X"21",  -- 33
        701 => X"22",  -- 34
        702 => X"23",  -- 35
        703 => X"24",  -- 36
        704 => X"26",  -- 38
        705 => X"28",  -- 40
        706 => X"2B",  -- 43
        707 => X"2D",  -- 45
        708 => X"2E",  -- 46
        709 => X"30",  -- 48
        710 => X"34",  -- 52
        711 => X"36",  -- 54
        712 => X"38",  -- 56
        713 => X"3A",  -- 58
        714 => X"3C",  -- 60
        715 => X"3E",  -- 62
        716 => X"3F",  -- 63
        717 => X"40",  -- 64
        718 => X"40",  -- 64
        719 => X"3F",  -- 63
        720 => X"41",  -- 65
        721 => X"42",  -- 66
        722 => X"41",  -- 65
        723 => X"42",  -- 66
        724 => X"42",  -- 66
        725 => X"42",  -- 66
        726 => X"42",  -- 66
        727 => X"42",  -- 66
        728 => X"40",  -- 64
        729 => X"40",  -- 64
        730 => X"44",  -- 68
        731 => X"50",  -- 80
        732 => X"61",  -- 97
        733 => X"70",  -- 112
        734 => X"78",  -- 120
        735 => X"7A",  -- 122
        736 => X"77",  -- 119
        737 => X"79",  -- 121
        738 => X"76",  -- 118
        739 => X"73",  -- 115
        740 => X"77",  -- 119
        741 => X"7C",  -- 124
        742 => X"77",  -- 119
        743 => X"6E",  -- 110
        744 => X"6E",  -- 110
        745 => X"54",  -- 84
        746 => X"45",  -- 69
        747 => X"53",  -- 83
        748 => X"59",  -- 89
        749 => X"42",  -- 66
        750 => X"2B",  -- 43
        751 => X"2F",  -- 47
        752 => X"3A",  -- 58
        753 => X"58",  -- 88
        754 => X"65",  -- 101
        755 => X"6A",  -- 106
        756 => X"76",  -- 118
        757 => X"75",  -- 117
        758 => X"6E",  -- 110
        759 => X"6F",  -- 111
        760 => X"79",  -- 121
        761 => X"65",  -- 101
        762 => X"55",  -- 85
        763 => X"44",  -- 68
        764 => X"2F",  -- 47
        765 => X"30",  -- 48
        766 => X"3B",  -- 59
        767 => X"39",  -- 57
        768 => X"3A",  -- 58
        769 => X"5F",  -- 95
        770 => X"78",  -- 120
        771 => X"89",  -- 137
        772 => X"88",  -- 136
        773 => X"88",  -- 136
        774 => X"9F",  -- 159
        775 => X"A7",  -- 167
        776 => X"A5",  -- 165
        777 => X"A4",  -- 164
        778 => X"A4",  -- 164
        779 => X"A5",  -- 165
        780 => X"A6",  -- 166
        781 => X"A7",  -- 167
        782 => X"A4",  -- 164
        783 => X"A4",  -- 164
        784 => X"A3",  -- 163
        785 => X"A1",  -- 161
        786 => X"A8",  -- 168
        787 => X"AA",  -- 170
        788 => X"A3",  -- 163
        789 => X"A3",  -- 163
        790 => X"A5",  -- 165
        791 => X"9F",  -- 159
        792 => X"9F",  -- 159
        793 => X"A0",  -- 160
        794 => X"A0",  -- 160
        795 => X"93",  -- 147
        796 => X"7B",  -- 123
        797 => X"6F",  -- 111
        798 => X"6D",  -- 109
        799 => X"65",  -- 101
        800 => X"51",  -- 81
        801 => X"52",  -- 82
        802 => X"4C",  -- 76
        803 => X"45",  -- 69
        804 => X"4E",  -- 78
        805 => X"61",  -- 97
        806 => X"6B",  -- 107
        807 => X"6B",  -- 107
        808 => X"79",  -- 121
        809 => X"7A",  -- 122
        810 => X"7A",  -- 122
        811 => X"7A",  -- 122
        812 => X"7B",  -- 123
        813 => X"7C",  -- 124
        814 => X"7F",  -- 127
        815 => X"82",  -- 130
        816 => X"85",  -- 133
        817 => X"86",  -- 134
        818 => X"86",  -- 134
        819 => X"84",  -- 132
        820 => X"86",  -- 134
        821 => X"87",  -- 135
        822 => X"8B",  -- 139
        823 => X"8E",  -- 142
        824 => X"8B",  -- 139
        825 => X"8C",  -- 140
        826 => X"91",  -- 145
        827 => X"94",  -- 148
        828 => X"90",  -- 144
        829 => X"88",  -- 136
        830 => X"88",  -- 136
        831 => X"8D",  -- 141
        832 => X"97",  -- 151
        833 => X"9A",  -- 154
        834 => X"9F",  -- 159
        835 => X"A1",  -- 161
        836 => X"A3",  -- 163
        837 => X"A6",  -- 166
        838 => X"AC",  -- 172
        839 => X"B0",  -- 176
        840 => X"AF",  -- 175
        841 => X"AD",  -- 173
        842 => X"AB",  -- 171
        843 => X"A9",  -- 169
        844 => X"A9",  -- 169
        845 => X"A9",  -- 169
        846 => X"A9",  -- 169
        847 => X"A8",  -- 168
        848 => X"AF",  -- 175
        849 => X"AD",  -- 173
        850 => X"AC",  -- 172
        851 => X"AE",  -- 174
        852 => X"B1",  -- 177
        853 => X"B5",  -- 181
        854 => X"B4",  -- 180
        855 => X"B3",  -- 179
        856 => X"AB",  -- 171
        857 => X"AC",  -- 172
        858 => X"AD",  -- 173
        859 => X"AC",  -- 172
        860 => X"AB",  -- 171
        861 => X"A8",  -- 168
        862 => X"A5",  -- 165
        863 => X"A3",  -- 163
        864 => X"99",  -- 153
        865 => X"97",  -- 151
        866 => X"97",  -- 151
        867 => X"9A",  -- 154
        868 => X"9B",  -- 155
        869 => X"99",  -- 153
        870 => X"96",  -- 150
        871 => X"96",  -- 150
        872 => X"9C",  -- 156
        873 => X"9C",  -- 156
        874 => X"9D",  -- 157
        875 => X"9E",  -- 158
        876 => X"9F",  -- 159
        877 => X"A0",  -- 160
        878 => X"9F",  -- 159
        879 => X"9D",  -- 157
        880 => X"A0",  -- 160
        881 => X"A2",  -- 162
        882 => X"A4",  -- 164
        883 => X"A6",  -- 166
        884 => X"A6",  -- 166
        885 => X"A8",  -- 168
        886 => X"AB",  -- 171
        887 => X"AD",  -- 173
        888 => X"AA",  -- 170
        889 => X"AB",  -- 171
        890 => X"AD",  -- 173
        891 => X"AD",  -- 173
        892 => X"AA",  -- 170
        893 => X"A0",  -- 160
        894 => X"94",  -- 148
        895 => X"8B",  -- 139
        896 => X"88",  -- 136
        897 => X"89",  -- 137
        898 => X"89",  -- 137
        899 => X"87",  -- 135
        900 => X"80",  -- 128
        901 => X"75",  -- 117
        902 => X"65",  -- 101
        903 => X"5A",  -- 90
        904 => X"4D",  -- 77
        905 => X"4E",  -- 78
        906 => X"4B",  -- 75
        907 => X"47",  -- 71
        908 => X"4D",  -- 77
        909 => X"58",  -- 88
        910 => X"5C",  -- 92
        911 => X"5C",  -- 92
        912 => X"5E",  -- 94
        913 => X"6C",  -- 108
        914 => X"78",  -- 120
        915 => X"86",  -- 134
        916 => X"99",  -- 153
        917 => X"A5",  -- 165
        918 => X"A8",  -- 168
        919 => X"AE",  -- 174
        920 => X"AC",  -- 172
        921 => X"AF",  -- 175
        922 => X"B3",  -- 179
        923 => X"B4",  -- 180
        924 => X"B3",  -- 179
        925 => X"B2",  -- 178
        926 => X"B4",  -- 180
        927 => X"B6",  -- 182
        928 => X"BD",  -- 189
        929 => X"BA",  -- 186
        930 => X"B9",  -- 185
        931 => X"BB",  -- 187
        932 => X"BE",  -- 190
        933 => X"BE",  -- 190
        934 => X"BA",  -- 186
        935 => X"B6",  -- 182
        936 => X"B5",  -- 181
        937 => X"B3",  -- 179
        938 => X"B2",  -- 178
        939 => X"B3",  -- 179
        940 => X"B6",  -- 182
        941 => X"B8",  -- 184
        942 => X"B7",  -- 183
        943 => X"B6",  -- 182
        944 => X"B5",  -- 181
        945 => X"B5",  -- 181
        946 => X"B5",  -- 181
        947 => X"B5",  -- 181
        948 => X"B5",  -- 181
        949 => X"B3",  -- 179
        950 => X"AF",  -- 175
        951 => X"AC",  -- 172
        952 => X"B5",  -- 181
        953 => X"B5",  -- 181
        954 => X"B8",  -- 184
        955 => X"BA",  -- 186
        956 => X"BA",  -- 186
        957 => X"B8",  -- 184
        958 => X"B2",  -- 178
        959 => X"AE",  -- 174
        960 => X"36",  -- 54
        961 => X"35",  -- 53
        962 => X"35",  -- 53
        963 => X"34",  -- 52
        964 => X"33",  -- 51
        965 => X"33",  -- 51
        966 => X"34",  -- 52
        967 => X"34",  -- 52
        968 => X"34",  -- 52
        969 => X"34",  -- 52
        970 => X"34",  -- 52
        971 => X"34",  -- 52
        972 => X"35",  -- 53
        973 => X"37",  -- 55
        974 => X"39",  -- 57
        975 => X"39",  -- 57
        976 => X"3A",  -- 58
        977 => X"3A",  -- 58
        978 => X"3A",  -- 58
        979 => X"3B",  -- 59
        980 => X"3B",  -- 59
        981 => X"3B",  -- 59
        982 => X"3B",  -- 59
        983 => X"3B",  -- 59
        984 => X"3B",  -- 59
        985 => X"3B",  -- 59
        986 => X"3C",  -- 60
        987 => X"3C",  -- 60
        988 => X"3C",  -- 60
        989 => X"3B",  -- 59
        990 => X"3A",  -- 58
        991 => X"3A",  -- 58
        992 => X"39",  -- 57
        993 => X"38",  -- 56
        994 => X"38",  -- 56
        995 => X"37",  -- 55
        996 => X"37",  -- 55
        997 => X"36",  -- 54
        998 => X"36",  -- 54
        999 => X"36",  -- 54
        1000 => X"34",  -- 52
        1001 => X"34",  -- 52
        1002 => X"32",  -- 50
        1003 => X"31",  -- 49
        1004 => X"30",  -- 48
        1005 => X"2F",  -- 47
        1006 => X"2E",  -- 46
        1007 => X"2E",  -- 46
        1008 => X"2D",  -- 45
        1009 => X"2C",  -- 44
        1010 => X"2C",  -- 44
        1011 => X"2B",  -- 43
        1012 => X"2A",  -- 42
        1013 => X"29",  -- 41
        1014 => X"29",  -- 41
        1015 => X"29",  -- 41
        1016 => X"25",  -- 37
        1017 => X"25",  -- 37
        1018 => X"24",  -- 36
        1019 => X"23",  -- 35
        1020 => X"24",  -- 36
        1021 => X"25",  -- 37
        1022 => X"26",  -- 38
        1023 => X"27",  -- 39
        1024 => X"2A",  -- 42
        1025 => X"2C",  -- 44
        1026 => X"2E",  -- 46
        1027 => X"30",  -- 48
        1028 => X"31",  -- 49
        1029 => X"33",  -- 51
        1030 => X"37",  -- 55
        1031 => X"39",  -- 57
        1032 => X"3B",  -- 59
        1033 => X"3D",  -- 61
        1034 => X"3F",  -- 63
        1035 => X"41",  -- 65
        1036 => X"43",  -- 67
        1037 => X"43",  -- 67
        1038 => X"43",  -- 67
        1039 => X"43",  -- 67
        1040 => X"44",  -- 68
        1041 => X"43",  -- 67
        1042 => X"44",  -- 68
        1043 => X"44",  -- 68
        1044 => X"43",  -- 67
        1045 => X"44",  -- 68
        1046 => X"43",  -- 67
        1047 => X"44",  -- 68
        1048 => X"45",  -- 69
        1049 => X"42",  -- 66
        1050 => X"44",  -- 68
        1051 => X"51",  -- 81
        1052 => X"65",  -- 101
        1053 => X"71",  -- 113
        1054 => X"72",  -- 114
        1055 => X"70",  -- 112
        1056 => X"6E",  -- 110
        1057 => X"6B",  -- 107
        1058 => X"62",  -- 98
        1059 => X"60",  -- 96
        1060 => X"66",  -- 102
        1061 => X"6E",  -- 110
        1062 => X"6E",  -- 110
        1063 => X"66",  -- 102
        1064 => X"6D",  -- 109
        1065 => X"57",  -- 87
        1066 => X"4B",  -- 75
        1067 => X"5C",  -- 92
        1068 => X"65",  -- 101
        1069 => X"45",  -- 69
        1070 => X"32",  -- 50
        1071 => X"44",  -- 68
        1072 => X"52",  -- 82
        1073 => X"63",  -- 99
        1074 => X"60",  -- 96
        1075 => X"62",  -- 98
        1076 => X"75",  -- 117
        1077 => X"72",  -- 114
        1078 => X"68",  -- 104
        1079 => X"76",  -- 118
        1080 => X"6C",  -- 108
        1081 => X"58",  -- 88
        1082 => X"4E",  -- 78
        1083 => X"3D",  -- 61
        1084 => X"25",  -- 37
        1085 => X"34",  -- 52
        1086 => X"4D",  -- 77
        1087 => X"46",  -- 70
        1088 => X"4E",  -- 78
        1089 => X"70",  -- 112
        1090 => X"87",  -- 135
        1091 => X"95",  -- 149
        1092 => X"91",  -- 145
        1093 => X"8F",  -- 143
        1094 => X"9F",  -- 159
        1095 => X"A3",  -- 163
        1096 => X"A4",  -- 164
        1097 => X"A3",  -- 163
        1098 => X"A4",  -- 164
        1099 => X"A4",  -- 164
        1100 => X"A5",  -- 165
        1101 => X"A5",  -- 165
        1102 => X"A4",  -- 164
        1103 => X"A1",  -- 161
        1104 => X"A4",  -- 164
        1105 => X"A5",  -- 165
        1106 => X"A8",  -- 168
        1107 => X"A8",  -- 168
        1108 => X"A3",  -- 163
        1109 => X"A1",  -- 161
        1110 => X"A3",  -- 163
        1111 => X"A4",  -- 164
        1112 => X"A8",  -- 168
        1113 => X"9F",  -- 159
        1114 => X"9A",  -- 154
        1115 => X"96",  -- 150
        1116 => X"91",  -- 145
        1117 => X"90",  -- 144
        1118 => X"87",  -- 135
        1119 => X"75",  -- 117
        1120 => X"68",  -- 104
        1121 => X"5F",  -- 95
        1122 => X"56",  -- 86
        1123 => X"5A",  -- 90
        1124 => X"6D",  -- 109
        1125 => X"79",  -- 121
        1126 => X"77",  -- 119
        1127 => X"6D",  -- 109
        1128 => X"7E",  -- 126
        1129 => X"7D",  -- 125
        1130 => X"7D",  -- 125
        1131 => X"7C",  -- 124
        1132 => X"7A",  -- 122
        1133 => X"7A",  -- 122
        1134 => X"7E",  -- 126
        1135 => X"81",  -- 129
        1136 => X"81",  -- 129
        1137 => X"82",  -- 130
        1138 => X"83",  -- 131
        1139 => X"83",  -- 131
        1140 => X"84",  -- 132
        1141 => X"88",  -- 136
        1142 => X"8C",  -- 140
        1143 => X"90",  -- 144
        1144 => X"8E",  -- 142
        1145 => X"8C",  -- 140
        1146 => X"8B",  -- 139
        1147 => X"8E",  -- 142
        1148 => X"90",  -- 144
        1149 => X"8E",  -- 142
        1150 => X"90",  -- 144
        1151 => X"96",  -- 150
        1152 => X"96",  -- 150
        1153 => X"97",  -- 151
        1154 => X"99",  -- 153
        1155 => X"9C",  -- 156
        1156 => X"A0",  -- 160
        1157 => X"A5",  -- 165
        1158 => X"AC",  -- 172
        1159 => X"B0",  -- 176
        1160 => X"AD",  -- 173
        1161 => X"AA",  -- 170
        1162 => X"A7",  -- 167
        1163 => X"A7",  -- 167
        1164 => X"AA",  -- 170
        1165 => X"AC",  -- 172
        1166 => X"AB",  -- 171
        1167 => X"AA",  -- 170
        1168 => X"B2",  -- 178
        1169 => X"B2",  -- 178
        1170 => X"B2",  -- 178
        1171 => X"B5",  -- 181
        1172 => X"B8",  -- 184
        1173 => X"BA",  -- 186
        1174 => X"B9",  -- 185
        1175 => X"B8",  -- 184
        1176 => X"B4",  -- 180
        1177 => X"B2",  -- 178
        1178 => X"B1",  -- 177
        1179 => X"B0",  -- 176
        1180 => X"B0",  -- 176
        1181 => X"AD",  -- 173
        1182 => X"A7",  -- 167
        1183 => X"A2",  -- 162
        1184 => X"A0",  -- 160
        1185 => X"9C",  -- 156
        1186 => X"98",  -- 152
        1187 => X"96",  -- 150
        1188 => X"97",  -- 151
        1189 => X"99",  -- 153
        1190 => X"9B",  -- 155
        1191 => X"9C",  -- 156
        1192 => X"9C",  -- 156
        1193 => X"9D",  -- 157
        1194 => X"A0",  -- 160
        1195 => X"A2",  -- 162
        1196 => X"A3",  -- 163
        1197 => X"A4",  -- 164
        1198 => X"A3",  -- 163
        1199 => X"A2",  -- 162
        1200 => X"A3",  -- 163
        1201 => X"A5",  -- 165
        1202 => X"A6",  -- 166
        1203 => X"A7",  -- 167
        1204 => X"A7",  -- 167
        1205 => X"A8",  -- 168
        1206 => X"AB",  -- 171
        1207 => X"AC",  -- 172
        1208 => X"AD",  -- 173
        1209 => X"AB",  -- 171
        1210 => X"AB",  -- 171
        1211 => X"AD",  -- 173
        1212 => X"AD",  -- 173
        1213 => X"A7",  -- 167
        1214 => X"9B",  -- 155
        1215 => X"90",  -- 144
        1216 => X"8B",  -- 139
        1217 => X"88",  -- 136
        1218 => X"87",  -- 135
        1219 => X"88",  -- 136
        1220 => X"88",  -- 136
        1221 => X"7E",  -- 126
        1222 => X"6D",  -- 109
        1223 => X"5F",  -- 95
        1224 => X"54",  -- 84
        1225 => X"56",  -- 86
        1226 => X"53",  -- 83
        1227 => X"4E",  -- 78
        1228 => X"4F",  -- 79
        1229 => X"55",  -- 85
        1230 => X"51",  -- 81
        1231 => X"49",  -- 73
        1232 => X"54",  -- 84
        1233 => X"61",  -- 97
        1234 => X"6A",  -- 106
        1235 => X"78",  -- 120
        1236 => X"8E",  -- 142
        1237 => X"9C",  -- 156
        1238 => X"A3",  -- 163
        1239 => X"AD",  -- 173
        1240 => X"AD",  -- 173
        1241 => X"B0",  -- 176
        1242 => X"B2",  -- 178
        1243 => X"B3",  -- 179
        1244 => X"B1",  -- 177
        1245 => X"B3",  -- 179
        1246 => X"B8",  -- 184
        1247 => X"BD",  -- 189
        1248 => X"BC",  -- 188
        1249 => X"BB",  -- 187
        1250 => X"BA",  -- 186
        1251 => X"BB",  -- 187
        1252 => X"BD",  -- 189
        1253 => X"BD",  -- 189
        1254 => X"B9",  -- 185
        1255 => X"B5",  -- 181
        1256 => X"B5",  -- 181
        1257 => X"B1",  -- 177
        1258 => X"AF",  -- 175
        1259 => X"B3",  -- 179
        1260 => X"B7",  -- 183
        1261 => X"BB",  -- 187
        1262 => X"B8",  -- 184
        1263 => X"B6",  -- 182
        1264 => X"B4",  -- 180
        1265 => X"B5",  -- 181
        1266 => X"B4",  -- 180
        1267 => X"B4",  -- 180
        1268 => X"B4",  -- 180
        1269 => X"B3",  -- 179
        1270 => X"AF",  -- 175
        1271 => X"AC",  -- 172
        1272 => X"B5",  -- 181
        1273 => X"B5",  -- 181
        1274 => X"B9",  -- 185
        1275 => X"BB",  -- 187
        1276 => X"BC",  -- 188
        1277 => X"BB",  -- 187
        1278 => X"B6",  -- 182
        1279 => X"B2",  -- 178
        1280 => X"37",  -- 55
        1281 => X"37",  -- 55
        1282 => X"36",  -- 54
        1283 => X"35",  -- 53
        1284 => X"34",  -- 52
        1285 => X"34",  -- 52
        1286 => X"34",  -- 52
        1287 => X"34",  -- 52
        1288 => X"35",  -- 53
        1289 => X"35",  -- 53
        1290 => X"35",  -- 53
        1291 => X"35",  -- 53
        1292 => X"36",  -- 54
        1293 => X"37",  -- 55
        1294 => X"39",  -- 57
        1295 => X"3A",  -- 58
        1296 => X"39",  -- 57
        1297 => X"39",  -- 57
        1298 => X"39",  -- 57
        1299 => X"3A",  -- 58
        1300 => X"3A",  -- 58
        1301 => X"3A",  -- 58
        1302 => X"3A",  -- 58
        1303 => X"3B",  -- 59
        1304 => X"3B",  -- 59
        1305 => X"3B",  -- 59
        1306 => X"3C",  -- 60
        1307 => X"3C",  -- 60
        1308 => X"3C",  -- 60
        1309 => X"3B",  -- 59
        1310 => X"3A",  -- 58
        1311 => X"3A",  -- 58
        1312 => X"39",  -- 57
        1313 => X"38",  -- 56
        1314 => X"38",  -- 56
        1315 => X"37",  -- 55
        1316 => X"37",  -- 55
        1317 => X"36",  -- 54
        1318 => X"36",  -- 54
        1319 => X"35",  -- 53
        1320 => X"34",  -- 52
        1321 => X"34",  -- 52
        1322 => X"32",  -- 50
        1323 => X"31",  -- 49
        1324 => X"30",  -- 48
        1325 => X"2F",  -- 47
        1326 => X"2E",  -- 46
        1327 => X"2E",  -- 46
        1328 => X"2D",  -- 45
        1329 => X"2C",  -- 44
        1330 => X"2C",  -- 44
        1331 => X"2B",  -- 43
        1332 => X"2A",  -- 42
        1333 => X"29",  -- 41
        1334 => X"29",  -- 41
        1335 => X"28",  -- 40
        1336 => X"25",  -- 37
        1337 => X"24",  -- 36
        1338 => X"23",  -- 35
        1339 => X"22",  -- 34
        1340 => X"23",  -- 35
        1341 => X"24",  -- 36
        1342 => X"25",  -- 37
        1343 => X"26",  -- 38
        1344 => X"29",  -- 41
        1345 => X"2B",  -- 43
        1346 => X"2E",  -- 46
        1347 => X"30",  -- 48
        1348 => X"31",  -- 49
        1349 => X"33",  -- 51
        1350 => X"36",  -- 54
        1351 => X"38",  -- 56
        1352 => X"3A",  -- 58
        1353 => X"3C",  -- 60
        1354 => X"3E",  -- 62
        1355 => X"41",  -- 65
        1356 => X"42",  -- 66
        1357 => X"43",  -- 67
        1358 => X"43",  -- 67
        1359 => X"43",  -- 67
        1360 => X"42",  -- 66
        1361 => X"42",  -- 66
        1362 => X"43",  -- 67
        1363 => X"42",  -- 66
        1364 => X"42",  -- 66
        1365 => X"43",  -- 67
        1366 => X"43",  -- 67
        1367 => X"43",  -- 67
        1368 => X"48",  -- 72
        1369 => X"42",  -- 66
        1370 => X"42",  -- 66
        1371 => X"4D",  -- 77
        1372 => X"61",  -- 97
        1373 => X"6A",  -- 106
        1374 => X"65",  -- 101
        1375 => X"5D",  -- 93
        1376 => X"5E",  -- 94
        1377 => X"57",  -- 87
        1378 => X"4C",  -- 76
        1379 => X"49",  -- 73
        1380 => X"4E",  -- 78
        1381 => X"59",  -- 89
        1382 => X"60",  -- 96
        1383 => X"60",  -- 96
        1384 => X"62",  -- 98
        1385 => X"57",  -- 87
        1386 => X"54",  -- 84
        1387 => X"67",  -- 103
        1388 => X"6C",  -- 108
        1389 => X"4A",  -- 74
        1390 => X"3C",  -- 60
        1391 => X"56",  -- 86
        1392 => X"64",  -- 100
        1393 => X"62",  -- 98
        1394 => X"51",  -- 81
        1395 => X"53",  -- 83
        1396 => X"6A",  -- 106
        1397 => X"69",  -- 105
        1398 => X"62",  -- 98
        1399 => X"72",  -- 114
        1400 => X"58",  -- 88
        1401 => X"46",  -- 70
        1402 => X"41",  -- 65
        1403 => X"36",  -- 54
        1404 => X"29",  -- 41
        1405 => X"45",  -- 69
        1406 => X"63",  -- 99
        1407 => X"5F",  -- 95
        1408 => X"67",  -- 103
        1409 => X"82",  -- 130
        1410 => X"8F",  -- 143
        1411 => X"97",  -- 151
        1412 => X"96",  -- 150
        1413 => X"96",  -- 150
        1414 => X"A1",  -- 161
        1415 => X"9B",  -- 155
        1416 => X"9F",  -- 159
        1417 => X"9E",  -- 158
        1418 => X"9E",  -- 158
        1419 => X"9F",  -- 159
        1420 => X"A1",  -- 161
        1421 => X"A1",  -- 161
        1422 => X"9F",  -- 159
        1423 => X"9F",  -- 159
        1424 => X"9D",  -- 157
        1425 => X"A1",  -- 161
        1426 => X"A1",  -- 161
        1427 => X"9D",  -- 157
        1428 => X"9D",  -- 157
        1429 => X"9D",  -- 157
        1430 => X"A0",  -- 160
        1431 => X"A5",  -- 165
        1432 => X"AD",  -- 173
        1433 => X"A1",  -- 161
        1434 => X"9B",  -- 155
        1435 => X"9C",  -- 156
        1436 => X"9D",  -- 157
        1437 => X"9D",  -- 157
        1438 => X"8F",  -- 143
        1439 => X"77",  -- 119
        1440 => X"73",  -- 115
        1441 => X"65",  -- 101
        1442 => X"64",  -- 100
        1443 => X"73",  -- 115
        1444 => X"7D",  -- 125
        1445 => X"7A",  -- 122
        1446 => X"73",  -- 115
        1447 => X"71",  -- 113
        1448 => X"76",  -- 118
        1449 => X"78",  -- 120
        1450 => X"7A",  -- 122
        1451 => X"7A",  -- 122
        1452 => X"7A",  -- 122
        1453 => X"7C",  -- 124
        1454 => X"81",  -- 129
        1455 => X"86",  -- 134
        1456 => X"7E",  -- 126
        1457 => X"7F",  -- 127
        1458 => X"82",  -- 130
        1459 => X"83",  -- 131
        1460 => X"85",  -- 133
        1461 => X"87",  -- 135
        1462 => X"8B",  -- 139
        1463 => X"8E",  -- 142
        1464 => X"8F",  -- 143
        1465 => X"8A",  -- 138
        1466 => X"88",  -- 136
        1467 => X"8A",  -- 138
        1468 => X"8E",  -- 142
        1469 => X"8F",  -- 143
        1470 => X"93",  -- 147
        1471 => X"95",  -- 149
        1472 => X"95",  -- 149
        1473 => X"94",  -- 148
        1474 => X"95",  -- 149
        1475 => X"98",  -- 152
        1476 => X"9D",  -- 157
        1477 => X"A3",  -- 163
        1478 => X"A6",  -- 166
        1479 => X"A8",  -- 168
        1480 => X"A9",  -- 169
        1481 => X"A7",  -- 167
        1482 => X"A5",  -- 165
        1483 => X"A7",  -- 167
        1484 => X"AB",  -- 171
        1485 => X"AE",  -- 174
        1486 => X"AF",  -- 175
        1487 => X"AE",  -- 174
        1488 => X"AD",  -- 173
        1489 => X"AF",  -- 175
        1490 => X"B2",  -- 178
        1491 => X"B6",  -- 182
        1492 => X"B7",  -- 183
        1493 => X"B8",  -- 184
        1494 => X"B6",  -- 182
        1495 => X"B4",  -- 180
        1496 => X"B5",  -- 181
        1497 => X"B2",  -- 178
        1498 => X"B0",  -- 176
        1499 => X"AE",  -- 174
        1500 => X"AE",  -- 174
        1501 => X"AB",  -- 171
        1502 => X"A5",  -- 165
        1503 => X"9F",  -- 159
        1504 => X"9E",  -- 158
        1505 => X"9B",  -- 155
        1506 => X"97",  -- 151
        1507 => X"94",  -- 148
        1508 => X"95",  -- 149
        1509 => X"99",  -- 153
        1510 => X"9B",  -- 155
        1511 => X"9C",  -- 156
        1512 => X"9C",  -- 156
        1513 => X"9E",  -- 158
        1514 => X"A1",  -- 161
        1515 => X"A3",  -- 163
        1516 => X"A5",  -- 165
        1517 => X"A6",  -- 166
        1518 => X"A7",  -- 167
        1519 => X"A7",  -- 167
        1520 => X"A3",  -- 163
        1521 => X"A4",  -- 164
        1522 => X"A5",  -- 165
        1523 => X"A5",  -- 165
        1524 => X"A5",  -- 165
        1525 => X"A5",  -- 165
        1526 => X"A7",  -- 167
        1527 => X"A8",  -- 168
        1528 => X"AF",  -- 175
        1529 => X"AB",  -- 171
        1530 => X"A9",  -- 169
        1531 => X"AA",  -- 170
        1532 => X"AE",  -- 174
        1533 => X"AB",  -- 171
        1534 => X"A2",  -- 162
        1535 => X"99",  -- 153
        1536 => X"8F",  -- 143
        1537 => X"89",  -- 137
        1538 => X"87",  -- 135
        1539 => X"8A",  -- 138
        1540 => X"8D",  -- 141
        1541 => X"88",  -- 136
        1542 => X"79",  -- 121
        1543 => X"6C",  -- 108
        1544 => X"64",  -- 100
        1545 => X"65",  -- 101
        1546 => X"5F",  -- 95
        1547 => X"53",  -- 83
        1548 => X"49",  -- 73
        1549 => X"46",  -- 70
        1550 => X"41",  -- 65
        1551 => X"3A",  -- 58
        1552 => X"50",  -- 80
        1553 => X"59",  -- 89
        1554 => X"5E",  -- 94
        1555 => X"66",  -- 102
        1556 => X"75",  -- 117
        1557 => X"82",  -- 130
        1558 => X"8D",  -- 141
        1559 => X"9C",  -- 156
        1560 => X"A2",  -- 162
        1561 => X"A9",  -- 169
        1562 => X"AF",  -- 175
        1563 => X"B2",  -- 178
        1564 => X"B2",  -- 178
        1565 => X"B4",  -- 180
        1566 => X"B8",  -- 184
        1567 => X"BD",  -- 189
        1568 => X"BB",  -- 187
        1569 => X"BB",  -- 187
        1570 => X"BB",  -- 187
        1571 => X"BC",  -- 188
        1572 => X"BB",  -- 187
        1573 => X"B9",  -- 185
        1574 => X"B6",  -- 182
        1575 => X"B6",  -- 182
        1576 => X"BD",  -- 189
        1577 => X"BA",  -- 186
        1578 => X"B6",  -- 182
        1579 => X"B5",  -- 181
        1580 => X"B7",  -- 183
        1581 => X"B6",  -- 182
        1582 => X"B2",  -- 178
        1583 => X"AD",  -- 173
        1584 => X"B4",  -- 180
        1585 => X"B3",  -- 179
        1586 => X"B2",  -- 178
        1587 => X"B2",  -- 178
        1588 => X"B2",  -- 178
        1589 => X"B2",  -- 178
        1590 => X"B1",  -- 177
        1591 => X"B0",  -- 176
        1592 => X"B5",  -- 181
        1593 => X"B5",  -- 181
        1594 => X"B9",  -- 185
        1595 => X"BB",  -- 187
        1596 => X"BD",  -- 189
        1597 => X"BE",  -- 190
        1598 => X"B9",  -- 185
        1599 => X"B6",  -- 182
        1600 => X"39",  -- 57
        1601 => X"38",  -- 56
        1602 => X"37",  -- 55
        1603 => X"36",  -- 54
        1604 => X"35",  -- 53
        1605 => X"35",  -- 53
        1606 => X"35",  -- 53
        1607 => X"35",  -- 53
        1608 => X"36",  -- 54
        1609 => X"36",  -- 54
        1610 => X"36",  -- 54
        1611 => X"36",  -- 54
        1612 => X"36",  -- 54
        1613 => X"37",  -- 55
        1614 => X"39",  -- 57
        1615 => X"3A",  -- 58
        1616 => X"39",  -- 57
        1617 => X"39",  -- 57
        1618 => X"39",  -- 57
        1619 => X"3A",  -- 58
        1620 => X"3A",  -- 58
        1621 => X"3A",  -- 58
        1622 => X"3A",  -- 58
        1623 => X"3A",  -- 58
        1624 => X"3B",  -- 59
        1625 => X"3B",  -- 59
        1626 => X"3C",  -- 60
        1627 => X"3C",  -- 60
        1628 => X"3C",  -- 60
        1629 => X"3B",  -- 59
        1630 => X"3A",  -- 58
        1631 => X"3A",  -- 58
        1632 => X"39",  -- 57
        1633 => X"38",  -- 56
        1634 => X"38",  -- 56
        1635 => X"37",  -- 55
        1636 => X"37",  -- 55
        1637 => X"36",  -- 54
        1638 => X"36",  -- 54
        1639 => X"35",  -- 53
        1640 => X"34",  -- 52
        1641 => X"34",  -- 52
        1642 => X"32",  -- 50
        1643 => X"31",  -- 49
        1644 => X"30",  -- 48
        1645 => X"2F",  -- 47
        1646 => X"2E",  -- 46
        1647 => X"2E",  -- 46
        1648 => X"2D",  -- 45
        1649 => X"2C",  -- 44
        1650 => X"2C",  -- 44
        1651 => X"2B",  -- 43
        1652 => X"2A",  -- 42
        1653 => X"29",  -- 41
        1654 => X"29",  -- 41
        1655 => X"28",  -- 40
        1656 => X"25",  -- 37
        1657 => X"24",  -- 36
        1658 => X"23",  -- 35
        1659 => X"22",  -- 34
        1660 => X"23",  -- 35
        1661 => X"24",  -- 36
        1662 => X"25",  -- 37
        1663 => X"26",  -- 38
        1664 => X"29",  -- 41
        1665 => X"2B",  -- 43
        1666 => X"2E",  -- 46
        1667 => X"2F",  -- 47
        1668 => X"31",  -- 49
        1669 => X"33",  -- 51
        1670 => X"36",  -- 54
        1671 => X"38",  -- 56
        1672 => X"3A",  -- 58
        1673 => X"3B",  -- 59
        1674 => X"3E",  -- 62
        1675 => X"40",  -- 64
        1676 => X"42",  -- 66
        1677 => X"43",  -- 67
        1678 => X"43",  -- 67
        1679 => X"43",  -- 67
        1680 => X"41",  -- 65
        1681 => X"41",  -- 65
        1682 => X"42",  -- 66
        1683 => X"42",  -- 66
        1684 => X"42",  -- 66
        1685 => X"42",  -- 66
        1686 => X"42",  -- 66
        1687 => X"42",  -- 66
        1688 => X"46",  -- 70
        1689 => X"41",  -- 65
        1690 => X"43",  -- 67
        1691 => X"4D",  -- 77
        1692 => X"59",  -- 89
        1693 => X"5A",  -- 90
        1694 => X"51",  -- 81
        1695 => X"46",  -- 70
        1696 => X"48",  -- 72
        1697 => X"43",  -- 67
        1698 => X"3D",  -- 61
        1699 => X"39",  -- 57
        1700 => X"3D",  -- 61
        1701 => X"47",  -- 71
        1702 => X"55",  -- 85
        1703 => X"5C",  -- 92
        1704 => X"5B",  -- 91
        1705 => X"5A",  -- 90
        1706 => X"65",  -- 101
        1707 => X"78",  -- 120
        1708 => X"75",  -- 117
        1709 => X"58",  -- 88
        1710 => X"50",  -- 80
        1711 => X"62",  -- 98
        1712 => X"69",  -- 105
        1713 => X"56",  -- 86
        1714 => X"40",  -- 64
        1715 => X"47",  -- 71
        1716 => X"5D",  -- 93
        1717 => X"5A",  -- 90
        1718 => X"55",  -- 85
        1719 => X"64",  -- 100
        1720 => X"47",  -- 71
        1721 => X"39",  -- 57
        1722 => X"36",  -- 54
        1723 => X"35",  -- 53
        1724 => X"3C",  -- 60
        1725 => X"59",  -- 89
        1726 => X"74",  -- 116
        1727 => X"73",  -- 115
        1728 => X"79",  -- 121
        1729 => X"8E",  -- 142
        1730 => X"92",  -- 146
        1731 => X"97",  -- 151
        1732 => X"97",  -- 151
        1733 => X"9A",  -- 154
        1734 => X"A0",  -- 160
        1735 => X"96",  -- 150
        1736 => X"9C",  -- 156
        1737 => X"9D",  -- 157
        1738 => X"9C",  -- 156
        1739 => X"9D",  -- 157
        1740 => X"9E",  -- 158
        1741 => X"9E",  -- 158
        1742 => X"9D",  -- 157
        1743 => X"9B",  -- 155
        1744 => X"95",  -- 149
        1745 => X"9C",  -- 156
        1746 => X"97",  -- 151
        1747 => X"96",  -- 150
        1748 => X"9D",  -- 157
        1749 => X"9F",  -- 159
        1750 => X"A0",  -- 160
        1751 => X"A8",  -- 168
        1752 => X"A2",  -- 162
        1753 => X"A2",  -- 162
        1754 => X"A7",  -- 167
        1755 => X"A7",  -- 167
        1756 => X"A0",  -- 160
        1757 => X"9E",  -- 158
        1758 => X"97",  -- 151
        1759 => X"89",  -- 137
        1760 => X"81",  -- 129
        1761 => X"7E",  -- 126
        1762 => X"86",  -- 134
        1763 => X"92",  -- 146
        1764 => X"8A",  -- 138
        1765 => X"76",  -- 118
        1766 => X"71",  -- 113
        1767 => X"7A",  -- 122
        1768 => X"74",  -- 116
        1769 => X"77",  -- 119
        1770 => X"7A",  -- 122
        1771 => X"79",  -- 121
        1772 => X"78",  -- 120
        1773 => X"79",  -- 121
        1774 => X"7B",  -- 123
        1775 => X"81",  -- 129
        1776 => X"7E",  -- 126
        1777 => X"80",  -- 128
        1778 => X"82",  -- 130
        1779 => X"84",  -- 132
        1780 => X"84",  -- 132
        1781 => X"86",  -- 134
        1782 => X"88",  -- 136
        1783 => X"89",  -- 137
        1784 => X"8B",  -- 139
        1785 => X"8A",  -- 138
        1786 => X"8B",  -- 139
        1787 => X"8E",  -- 142
        1788 => X"90",  -- 144
        1789 => X"92",  -- 146
        1790 => X"92",  -- 146
        1791 => X"92",  -- 146
        1792 => X"97",  -- 151
        1793 => X"96",  -- 150
        1794 => X"95",  -- 149
        1795 => X"98",  -- 152
        1796 => X"9D",  -- 157
        1797 => X"A1",  -- 161
        1798 => X"A1",  -- 161
        1799 => X"A0",  -- 160
        1800 => X"A3",  -- 163
        1801 => X"A4",  -- 164
        1802 => X"A6",  -- 166
        1803 => X"A8",  -- 168
        1804 => X"AC",  -- 172
        1805 => X"AF",  -- 175
        1806 => X"B0",  -- 176
        1807 => X"B0",  -- 176
        1808 => X"AA",  -- 170
        1809 => X"AC",  -- 172
        1810 => X"B0",  -- 176
        1811 => X"B4",  -- 180
        1812 => X"B4",  -- 180
        1813 => X"B5",  -- 181
        1814 => X"B2",  -- 178
        1815 => X"B1",  -- 177
        1816 => X"B4",  -- 180
        1817 => X"B1",  -- 177
        1818 => X"AE",  -- 174
        1819 => X"AC",  -- 172
        1820 => X"AC",  -- 172
        1821 => X"AA",  -- 170
        1822 => X"A7",  -- 167
        1823 => X"A2",  -- 162
        1824 => X"98",  -- 152
        1825 => X"99",  -- 153
        1826 => X"99",  -- 153
        1827 => X"98",  -- 152
        1828 => X"9A",  -- 154
        1829 => X"9C",  -- 156
        1830 => X"9B",  -- 155
        1831 => X"98",  -- 152
        1832 => X"9B",  -- 155
        1833 => X"9E",  -- 158
        1834 => X"A0",  -- 160
        1835 => X"A2",  -- 162
        1836 => X"A2",  -- 162
        1837 => X"A3",  -- 163
        1838 => X"A5",  -- 165
        1839 => X"A7",  -- 167
        1840 => X"A4",  -- 164
        1841 => X"A5",  -- 165
        1842 => X"A7",  -- 167
        1843 => X"A7",  -- 167
        1844 => X"A7",  -- 167
        1845 => X"A6",  -- 166
        1846 => X"A8",  -- 168
        1847 => X"AA",  -- 170
        1848 => X"AE",  -- 174
        1849 => X"AA",  -- 170
        1850 => X"A8",  -- 168
        1851 => X"AA",  -- 170
        1852 => X"AE",  -- 174
        1853 => X"AD",  -- 173
        1854 => X"A7",  -- 167
        1855 => X"A0",  -- 160
        1856 => X"93",  -- 147
        1857 => X"8E",  -- 142
        1858 => X"8A",  -- 138
        1859 => X"8A",  -- 138
        1860 => X"8E",  -- 142
        1861 => X"8C",  -- 140
        1862 => X"84",  -- 132
        1863 => X"79",  -- 121
        1864 => X"74",  -- 116
        1865 => X"71",  -- 113
        1866 => X"68",  -- 104
        1867 => X"5E",  -- 94
        1868 => X"52",  -- 82
        1869 => X"4A",  -- 74
        1870 => X"47",  -- 71
        1871 => X"49",  -- 73
        1872 => X"56",  -- 86
        1873 => X"5B",  -- 91
        1874 => X"58",  -- 88
        1875 => X"57",  -- 87
        1876 => X"60",  -- 96
        1877 => X"68",  -- 104
        1878 => X"74",  -- 116
        1879 => X"85",  -- 133
        1880 => X"8E",  -- 142
        1881 => X"98",  -- 152
        1882 => X"A7",  -- 167
        1883 => X"B0",  -- 176
        1884 => X"B3",  -- 179
        1885 => X"B6",  -- 182
        1886 => X"B7",  -- 183
        1887 => X"BB",  -- 187
        1888 => X"BE",  -- 190
        1889 => X"BF",  -- 191
        1890 => X"C1",  -- 193
        1891 => X"C0",  -- 192
        1892 => X"BE",  -- 190
        1893 => X"BA",  -- 186
        1894 => X"BA",  -- 186
        1895 => X"B9",  -- 185
        1896 => X"B8",  -- 184
        1897 => X"B6",  -- 182
        1898 => X"B5",  -- 181
        1899 => X"B6",  -- 182
        1900 => X"B7",  -- 183
        1901 => X"B5",  -- 181
        1902 => X"B2",  -- 178
        1903 => X"AE",  -- 174
        1904 => X"B3",  -- 179
        1905 => X"B2",  -- 178
        1906 => X"B0",  -- 176
        1907 => X"B0",  -- 176
        1908 => X"B0",  -- 176
        1909 => X"B0",  -- 176
        1910 => X"B0",  -- 176
        1911 => X"AF",  -- 175
        1912 => X"B2",  -- 178
        1913 => X"B3",  -- 179
        1914 => X"B6",  -- 182
        1915 => X"B9",  -- 185
        1916 => X"BB",  -- 187
        1917 => X"BB",  -- 187
        1918 => X"B8",  -- 184
        1919 => X"B6",  -- 182
        1920 => X"3B",  -- 59
        1921 => X"3B",  -- 59
        1922 => X"3A",  -- 58
        1923 => X"39",  -- 57
        1924 => X"37",  -- 55
        1925 => X"37",  -- 55
        1926 => X"37",  -- 55
        1927 => X"37",  -- 55
        1928 => X"38",  -- 56
        1929 => X"38",  -- 56
        1930 => X"38",  -- 56
        1931 => X"38",  -- 56
        1932 => X"38",  -- 56
        1933 => X"39",  -- 57
        1934 => X"3B",  -- 59
        1935 => X"3C",  -- 60
        1936 => X"3C",  -- 60
        1937 => X"3C",  -- 60
        1938 => X"3C",  -- 60
        1939 => X"3C",  -- 60
        1940 => X"3D",  -- 61
        1941 => X"3D",  -- 61
        1942 => X"3D",  -- 61
        1943 => X"3D",  -- 61
        1944 => X"3D",  -- 61
        1945 => X"3D",  -- 61
        1946 => X"3D",  -- 61
        1947 => X"3D",  -- 61
        1948 => X"3D",  -- 61
        1949 => X"3C",  -- 60
        1950 => X"3C",  -- 60
        1951 => X"3B",  -- 59
        1952 => X"3A",  -- 58
        1953 => X"3A",  -- 58
        1954 => X"39",  -- 57
        1955 => X"39",  -- 57
        1956 => X"39",  -- 57
        1957 => X"38",  -- 56
        1958 => X"37",  -- 55
        1959 => X"37",  -- 55
        1960 => X"36",  -- 54
        1961 => X"35",  -- 53
        1962 => X"34",  -- 52
        1963 => X"33",  -- 51
        1964 => X"32",  -- 50
        1965 => X"31",  -- 49
        1966 => X"30",  -- 48
        1967 => X"2F",  -- 47
        1968 => X"2E",  -- 46
        1969 => X"2E",  -- 46
        1970 => X"2D",  -- 45
        1971 => X"2D",  -- 45
        1972 => X"2C",  -- 44
        1973 => X"2B",  -- 43
        1974 => X"2A",  -- 42
        1975 => X"2A",  -- 42
        1976 => X"26",  -- 38
        1977 => X"26",  -- 38
        1978 => X"25",  -- 37
        1979 => X"24",  -- 36
        1980 => X"25",  -- 37
        1981 => X"26",  -- 38
        1982 => X"27",  -- 39
        1983 => X"28",  -- 40
        1984 => X"2A",  -- 42
        1985 => X"2C",  -- 44
        1986 => X"2F",  -- 47
        1987 => X"31",  -- 49
        1988 => X"32",  -- 50
        1989 => X"34",  -- 52
        1990 => X"37",  -- 55
        1991 => X"39",  -- 57
        1992 => X"3B",  -- 59
        1993 => X"3C",  -- 60
        1994 => X"3F",  -- 63
        1995 => X"41",  -- 65
        1996 => X"43",  -- 67
        1997 => X"45",  -- 69
        1998 => X"45",  -- 69
        1999 => X"45",  -- 69
        2000 => X"43",  -- 67
        2001 => X"43",  -- 67
        2002 => X"44",  -- 68
        2003 => X"44",  -- 68
        2004 => X"43",  -- 67
        2005 => X"43",  -- 67
        2006 => X"44",  -- 68
        2007 => X"44",  -- 68
        2008 => X"44",  -- 68
        2009 => X"49",  -- 73
        2010 => X"51",  -- 81
        2011 => X"57",  -- 87
        2012 => X"58",  -- 88
        2013 => X"4F",  -- 79
        2014 => X"44",  -- 68
        2015 => X"3B",  -- 59
        2016 => X"36",  -- 54
        2017 => X"3C",  -- 60
        2018 => X"3F",  -- 63
        2019 => X"41",  -- 65
        2020 => X"42",  -- 66
        2021 => X"4A",  -- 74
        2022 => X"57",  -- 87
        2023 => X"63",  -- 99
        2024 => X"63",  -- 99
        2025 => X"64",  -- 100
        2026 => X"75",  -- 117
        2027 => X"82",  -- 130
        2028 => X"7A",  -- 122
        2029 => X"6A",  -- 106
        2030 => X"69",  -- 105
        2031 => X"6E",  -- 110
        2032 => X"67",  -- 103
        2033 => X"4A",  -- 74
        2034 => X"3C",  -- 60
        2035 => X"49",  -- 73
        2036 => X"56",  -- 86
        2037 => X"4E",  -- 78
        2038 => X"4A",  -- 74
        2039 => X"53",  -- 83
        2040 => X"45",  -- 69
        2041 => X"3C",  -- 60
        2042 => X"37",  -- 55
        2043 => X"42",  -- 66
        2044 => X"59",  -- 89
        2045 => X"72",  -- 114
        2046 => X"81",  -- 129
        2047 => X"83",  -- 131
        2048 => X"87",  -- 135
        2049 => X"99",  -- 153
        2050 => X"98",  -- 152
        2051 => X"99",  -- 153
        2052 => X"98",  -- 152
        2053 => X"99",  -- 153
        2054 => X"9E",  -- 158
        2055 => X"91",  -- 145
        2056 => X"9C",  -- 156
        2057 => X"9A",  -- 154
        2058 => X"99",  -- 153
        2059 => X"99",  -- 153
        2060 => X"9B",  -- 155
        2061 => X"9A",  -- 154
        2062 => X"97",  -- 151
        2063 => X"96",  -- 150
        2064 => X"94",  -- 148
        2065 => X"9B",  -- 155
        2066 => X"97",  -- 151
        2067 => X"96",  -- 150
        2068 => X"A1",  -- 161
        2069 => X"A1",  -- 161
        2070 => X"9C",  -- 156
        2071 => X"A5",  -- 165
        2072 => X"9B",  -- 155
        2073 => X"A0",  -- 160
        2074 => X"AB",  -- 171
        2075 => X"AC",  -- 172
        2076 => X"A5",  -- 165
        2077 => X"A6",  -- 166
        2078 => X"A9",  -- 169
        2079 => X"A4",  -- 164
        2080 => X"9C",  -- 156
        2081 => X"9D",  -- 157
        2082 => X"A2",  -- 162
        2083 => X"A4",  -- 164
        2084 => X"95",  -- 149
        2085 => X"7D",  -- 125
        2086 => X"73",  -- 115
        2087 => X"77",  -- 119
        2088 => X"72",  -- 114
        2089 => X"77",  -- 119
        2090 => X"7A",  -- 122
        2091 => X"7A",  -- 122
        2092 => X"75",  -- 117
        2093 => X"72",  -- 114
        2094 => X"76",  -- 118
        2095 => X"79",  -- 121
        2096 => X"7E",  -- 126
        2097 => X"7F",  -- 127
        2098 => X"81",  -- 129
        2099 => X"81",  -- 129
        2100 => X"82",  -- 130
        2101 => X"85",  -- 133
        2102 => X"86",  -- 134
        2103 => X"8A",  -- 138
        2104 => X"8A",  -- 138
        2105 => X"8B",  -- 139
        2106 => X"8D",  -- 141
        2107 => X"8F",  -- 143
        2108 => X"92",  -- 146
        2109 => X"94",  -- 148
        2110 => X"94",  -- 148
        2111 => X"93",  -- 147
        2112 => X"99",  -- 153
        2113 => X"97",  -- 151
        2114 => X"98",  -- 152
        2115 => X"9C",  -- 156
        2116 => X"A2",  -- 162
        2117 => X"A4",  -- 164
        2118 => X"A1",  -- 161
        2119 => X"9E",  -- 158
        2120 => X"9D",  -- 157
        2121 => X"A0",  -- 160
        2122 => X"A5",  -- 165
        2123 => X"A8",  -- 168
        2124 => X"AA",  -- 170
        2125 => X"AB",  -- 171
        2126 => X"AD",  -- 173
        2127 => X"AE",  -- 174
        2128 => X"AD",  -- 173
        2129 => X"AF",  -- 175
        2130 => X"B0",  -- 176
        2131 => X"B2",  -- 178
        2132 => X"B1",  -- 177
        2133 => X"B3",  -- 179
        2134 => X"B3",  -- 179
        2135 => X"B3",  -- 179
        2136 => X"B6",  -- 182
        2137 => X"B3",  -- 179
        2138 => X"B1",  -- 177
        2139 => X"AC",  -- 172
        2140 => X"AB",  -- 171
        2141 => X"A8",  -- 168
        2142 => X"A6",  -- 166
        2143 => X"A4",  -- 164
        2144 => X"99",  -- 153
        2145 => X"9A",  -- 154
        2146 => X"9A",  -- 154
        2147 => X"97",  -- 151
        2148 => X"9A",  -- 154
        2149 => X"9E",  -- 158
        2150 => X"9E",  -- 158
        2151 => X"9B",  -- 155
        2152 => X"9D",  -- 157
        2153 => X"9E",  -- 158
        2154 => X"A0",  -- 160
        2155 => X"9F",  -- 159
        2156 => X"9E",  -- 158
        2157 => X"9E",  -- 158
        2158 => X"A0",  -- 160
        2159 => X"A3",  -- 163
        2160 => X"A5",  -- 165
        2161 => X"A7",  -- 167
        2162 => X"A9",  -- 169
        2163 => X"AA",  -- 170
        2164 => X"AA",  -- 170
        2165 => X"AB",  -- 171
        2166 => X"AD",  -- 173
        2167 => X"AE",  -- 174
        2168 => X"AD",  -- 173
        2169 => X"AC",  -- 172
        2170 => X"AC",  -- 172
        2171 => X"AF",  -- 175
        2172 => X"B3",  -- 179
        2173 => X"B1",  -- 177
        2174 => X"AC",  -- 172
        2175 => X"A7",  -- 167
        2176 => X"99",  -- 153
        2177 => X"95",  -- 149
        2178 => X"8F",  -- 143
        2179 => X"8C",  -- 140
        2180 => X"8E",  -- 142
        2181 => X"8E",  -- 142
        2182 => X"8B",  -- 139
        2183 => X"88",  -- 136
        2184 => X"82",  -- 130
        2185 => X"7B",  -- 123
        2186 => X"78",  -- 120
        2187 => X"77",  -- 119
        2188 => X"70",  -- 112
        2189 => X"63",  -- 99
        2190 => X"5D",  -- 93
        2191 => X"60",  -- 96
        2192 => X"63",  -- 99
        2193 => X"5E",  -- 94
        2194 => X"53",  -- 83
        2195 => X"50",  -- 80
        2196 => X"55",  -- 85
        2197 => X"58",  -- 88
        2198 => X"5C",  -- 92
        2199 => X"69",  -- 105
        2200 => X"75",  -- 117
        2201 => X"81",  -- 129
        2202 => X"93",  -- 147
        2203 => X"9E",  -- 158
        2204 => X"A4",  -- 164
        2205 => X"AA",  -- 170
        2206 => X"B4",  -- 180
        2207 => X"B9",  -- 185
        2208 => X"C1",  -- 193
        2209 => X"C0",  -- 192
        2210 => X"BE",  -- 190
        2211 => X"BE",  -- 190
        2212 => X"BE",  -- 190
        2213 => X"BD",  -- 189
        2214 => X"B9",  -- 185
        2215 => X"B6",  -- 182
        2216 => X"AC",  -- 172
        2217 => X"AF",  -- 175
        2218 => X"B2",  -- 178
        2219 => X"B6",  -- 182
        2220 => X"B9",  -- 185
        2221 => X"B9",  -- 185
        2222 => X"B8",  -- 184
        2223 => X"B7",  -- 183
        2224 => X"B5",  -- 181
        2225 => X"B3",  -- 179
        2226 => X"B3",  -- 179
        2227 => X"B3",  -- 179
        2228 => X"B1",  -- 177
        2229 => X"AF",  -- 175
        2230 => X"AD",  -- 173
        2231 => X"AA",  -- 170
        2232 => X"AC",  -- 172
        2233 => X"AC",  -- 172
        2234 => X"B0",  -- 176
        2235 => X"B2",  -- 178
        2236 => X"B5",  -- 181
        2237 => X"B5",  -- 181
        2238 => X"B3",  -- 179
        2239 => X"B1",  -- 177
        2240 => X"3B",  -- 59
        2241 => X"3A",  -- 58
        2242 => X"39",  -- 57
        2243 => X"38",  -- 56
        2244 => X"36",  -- 54
        2245 => X"36",  -- 54
        2246 => X"36",  -- 54
        2247 => X"36",  -- 54
        2248 => X"38",  -- 56
        2249 => X"38",  -- 56
        2250 => X"37",  -- 55
        2251 => X"37",  -- 55
        2252 => X"38",  -- 56
        2253 => X"38",  -- 56
        2254 => X"3A",  -- 58
        2255 => X"3B",  -- 59
        2256 => X"3C",  -- 60
        2257 => X"3C",  -- 60
        2258 => X"3C",  -- 60
        2259 => X"3C",  -- 60
        2260 => X"3D",  -- 61
        2261 => X"3D",  -- 61
        2262 => X"3D",  -- 61
        2263 => X"3D",  -- 61
        2264 => X"3C",  -- 60
        2265 => X"3C",  -- 60
        2266 => X"3C",  -- 60
        2267 => X"3C",  -- 60
        2268 => X"3C",  -- 60
        2269 => X"3B",  -- 59
        2270 => X"3B",  -- 59
        2271 => X"3A",  -- 58
        2272 => X"39",  -- 57
        2273 => X"39",  -- 57
        2274 => X"38",  -- 56
        2275 => X"37",  -- 55
        2276 => X"38",  -- 56
        2277 => X"37",  -- 55
        2278 => X"36",  -- 54
        2279 => X"36",  -- 54
        2280 => X"35",  -- 53
        2281 => X"34",  -- 52
        2282 => X"33",  -- 51
        2283 => X"32",  -- 50
        2284 => X"31",  -- 49
        2285 => X"2F",  -- 47
        2286 => X"2F",  -- 47
        2287 => X"2E",  -- 46
        2288 => X"2D",  -- 45
        2289 => X"2D",  -- 45
        2290 => X"2C",  -- 44
        2291 => X"2B",  -- 43
        2292 => X"2B",  -- 43
        2293 => X"2A",  -- 42
        2294 => X"29",  -- 41
        2295 => X"29",  -- 41
        2296 => X"26",  -- 38
        2297 => X"25",  -- 37
        2298 => X"24",  -- 36
        2299 => X"24",  -- 36
        2300 => X"24",  -- 36
        2301 => X"25",  -- 37
        2302 => X"26",  -- 38
        2303 => X"27",  -- 39
        2304 => X"29",  -- 41
        2305 => X"2B",  -- 43
        2306 => X"2E",  -- 46
        2307 => X"30",  -- 48
        2308 => X"31",  -- 49
        2309 => X"33",  -- 51
        2310 => X"36",  -- 54
        2311 => X"38",  -- 56
        2312 => X"39",  -- 57
        2313 => X"3B",  -- 59
        2314 => X"3D",  -- 61
        2315 => X"40",  -- 64
        2316 => X"42",  -- 66
        2317 => X"44",  -- 68
        2318 => X"44",  -- 68
        2319 => X"44",  -- 68
        2320 => X"43",  -- 67
        2321 => X"44",  -- 68
        2322 => X"44",  -- 68
        2323 => X"43",  -- 67
        2324 => X"44",  -- 68
        2325 => X"43",  -- 67
        2326 => X"44",  -- 68
        2327 => X"44",  -- 68
        2328 => X"47",  -- 71
        2329 => X"54",  -- 84
        2330 => X"62",  -- 98
        2331 => X"66",  -- 102
        2332 => X"5D",  -- 93
        2333 => X"4D",  -- 77
        2334 => X"40",  -- 64
        2335 => X"3A",  -- 58
        2336 => X"32",  -- 50
        2337 => X"3E",  -- 62
        2338 => X"4B",  -- 75
        2339 => X"51",  -- 81
        2340 => X"50",  -- 80
        2341 => X"54",  -- 84
        2342 => X"62",  -- 98
        2343 => X"6F",  -- 111
        2344 => X"6F",  -- 111
        2345 => X"6C",  -- 108
        2346 => X"7B",  -- 123
        2347 => X"81",  -- 129
        2348 => X"76",  -- 118
        2349 => X"73",  -- 115
        2350 => X"7B",  -- 123
        2351 => X"76",  -- 118
        2352 => X"60",  -- 96
        2353 => X"42",  -- 66
        2354 => X"3C",  -- 60
        2355 => X"4E",  -- 78
        2356 => X"52",  -- 82
        2357 => X"45",  -- 69
        2358 => X"42",  -- 66
        2359 => X"45",  -- 69
        2360 => X"4C",  -- 76
        2361 => X"45",  -- 69
        2362 => X"40",  -- 64
        2363 => X"50",  -- 80
        2364 => X"72",  -- 114
        2365 => X"85",  -- 133
        2366 => X"88",  -- 136
        2367 => X"8B",  -- 139
        2368 => X"90",  -- 144
        2369 => X"A2",  -- 162
        2370 => X"A1",  -- 161
        2371 => X"9D",  -- 157
        2372 => X"9A",  -- 154
        2373 => X"98",  -- 152
        2374 => X"9D",  -- 157
        2375 => X"8E",  -- 142
        2376 => X"97",  -- 151
        2377 => X"96",  -- 150
        2378 => X"94",  -- 148
        2379 => X"94",  -- 148
        2380 => X"92",  -- 146
        2381 => X"91",  -- 145
        2382 => X"90",  -- 144
        2383 => X"8E",  -- 142
        2384 => X"93",  -- 147
        2385 => X"9C",  -- 156
        2386 => X"95",  -- 149
        2387 => X"96",  -- 150
        2388 => X"A3",  -- 163
        2389 => X"9F",  -- 159
        2390 => X"95",  -- 149
        2391 => X"9B",  -- 155
        2392 => X"A0",  -- 160
        2393 => X"A2",  -- 162
        2394 => X"A7",  -- 167
        2395 => X"A8",  -- 168
        2396 => X"A5",  -- 165
        2397 => X"AA",  -- 170
        2398 => X"B1",  -- 177
        2399 => X"AB",  -- 171
        2400 => X"AF",  -- 175
        2401 => X"AC",  -- 172
        2402 => X"A7",  -- 167
        2403 => X"A0",  -- 160
        2404 => X"94",  -- 148
        2405 => X"83",  -- 131
        2406 => X"72",  -- 114
        2407 => X"65",  -- 101
        2408 => X"69",  -- 105
        2409 => X"6E",  -- 110
        2410 => X"75",  -- 117
        2411 => X"77",  -- 119
        2412 => X"75",  -- 117
        2413 => X"75",  -- 117
        2414 => X"78",  -- 120
        2415 => X"7C",  -- 124
        2416 => X"7B",  -- 123
        2417 => X"7C",  -- 124
        2418 => X"7E",  -- 126
        2419 => X"7F",  -- 127
        2420 => X"80",  -- 128
        2421 => X"84",  -- 132
        2422 => X"8A",  -- 138
        2423 => X"8D",  -- 141
        2424 => X"8A",  -- 138
        2425 => X"8D",  -- 141
        2426 => X"8D",  -- 141
        2427 => X"8C",  -- 140
        2428 => X"8E",  -- 142
        2429 => X"93",  -- 147
        2430 => X"97",  -- 151
        2431 => X"98",  -- 152
        2432 => X"98",  -- 152
        2433 => X"97",  -- 151
        2434 => X"99",  -- 153
        2435 => X"9F",  -- 159
        2436 => X"A6",  -- 166
        2437 => X"A9",  -- 169
        2438 => X"A5",  -- 165
        2439 => X"A1",  -- 161
        2440 => X"99",  -- 153
        2441 => X"9E",  -- 158
        2442 => X"A4",  -- 164
        2443 => X"A7",  -- 167
        2444 => X"A7",  -- 167
        2445 => X"A7",  -- 167
        2446 => X"A9",  -- 169
        2447 => X"AA",  -- 170
        2448 => X"B0",  -- 176
        2449 => X"AF",  -- 175
        2450 => X"AF",  -- 175
        2451 => X"AE",  -- 174
        2452 => X"AD",  -- 173
        2453 => X"B0",  -- 176
        2454 => X"B2",  -- 178
        2455 => X"B5",  -- 181
        2456 => X"B8",  -- 184
        2457 => X"B5",  -- 181
        2458 => X"B1",  -- 177
        2459 => X"AA",  -- 170
        2460 => X"A6",  -- 166
        2461 => X"A2",  -- 162
        2462 => X"A0",  -- 160
        2463 => X"9F",  -- 159
        2464 => X"9A",  -- 154
        2465 => X"9A",  -- 154
        2466 => X"95",  -- 149
        2467 => X"90",  -- 144
        2468 => X"92",  -- 146
        2469 => X"9A",  -- 154
        2470 => X"9F",  -- 159
        2471 => X"9F",  -- 159
        2472 => X"9F",  -- 159
        2473 => X"A0",  -- 160
        2474 => X"A0",  -- 160
        2475 => X"9E",  -- 158
        2476 => X"9B",  -- 155
        2477 => X"9B",  -- 155
        2478 => X"9D",  -- 157
        2479 => X"9F",  -- 159
        2480 => X"A2",  -- 162
        2481 => X"A4",  -- 164
        2482 => X"A7",  -- 167
        2483 => X"A9",  -- 169
        2484 => X"AA",  -- 170
        2485 => X"AC",  -- 172
        2486 => X"AE",  -- 174
        2487 => X"B0",  -- 176
        2488 => X"AD",  -- 173
        2489 => X"AE",  -- 174
        2490 => X"B1",  -- 177
        2491 => X"B5",  -- 181
        2492 => X"B8",  -- 184
        2493 => X"B6",  -- 182
        2494 => X"B0",  -- 176
        2495 => X"AB",  -- 171
        2496 => X"A1",  -- 161
        2497 => X"9C",  -- 156
        2498 => X"94",  -- 148
        2499 => X"90",  -- 144
        2500 => X"8F",  -- 143
        2501 => X"8F",  -- 143
        2502 => X"91",  -- 145
        2503 => X"92",  -- 146
        2504 => X"8F",  -- 143
        2505 => X"89",  -- 137
        2506 => X"89",  -- 137
        2507 => X"90",  -- 144
        2508 => X"89",  -- 137
        2509 => X"73",  -- 115
        2510 => X"64",  -- 100
        2511 => X"62",  -- 98
        2512 => X"67",  -- 103
        2513 => X"5F",  -- 95
        2514 => X"50",  -- 80
        2515 => X"4B",  -- 75
        2516 => X"50",  -- 80
        2517 => X"4E",  -- 78
        2518 => X"4B",  -- 75
        2519 => X"54",  -- 84
        2520 => X"62",  -- 98
        2521 => X"6B",  -- 107
        2522 => X"78",  -- 120
        2523 => X"82",  -- 130
        2524 => X"8C",  -- 140
        2525 => X"9A",  -- 154
        2526 => X"AA",  -- 170
        2527 => X"B6",  -- 182
        2528 => X"BE",  -- 190
        2529 => X"B9",  -- 185
        2530 => X"B4",  -- 180
        2531 => X"B6",  -- 182
        2532 => X"B9",  -- 185
        2533 => X"B9",  -- 185
        2534 => X"B4",  -- 180
        2535 => X"AC",  -- 172
        2536 => X"AD",  -- 173
        2537 => X"B1",  -- 177
        2538 => X"B5",  -- 181
        2539 => X"B9",  -- 185
        2540 => X"BA",  -- 186
        2541 => X"B9",  -- 185
        2542 => X"B8",  -- 184
        2543 => X"B7",  -- 183
        2544 => X"B8",  -- 184
        2545 => X"B7",  -- 183
        2546 => X"B8",  -- 184
        2547 => X"B7",  -- 183
        2548 => X"B4",  -- 180
        2549 => X"AF",  -- 175
        2550 => X"AA",  -- 170
        2551 => X"A5",  -- 165
        2552 => X"A7",  -- 167
        2553 => X"A8",  -- 168
        2554 => X"AA",  -- 170
        2555 => X"AC",  -- 172
        2556 => X"AF",  -- 175
        2557 => X"AF",  -- 175
        2558 => X"AD",  -- 173
        2559 => X"AB",  -- 171
        2560 => X"3D",  -- 61
        2561 => X"3C",  -- 60
        2562 => X"3A",  -- 58
        2563 => X"39",  -- 57
        2564 => X"37",  -- 55
        2565 => X"37",  -- 55
        2566 => X"38",  -- 56
        2567 => X"39",  -- 57
        2568 => X"39",  -- 57
        2569 => X"39",  -- 57
        2570 => X"39",  -- 57
        2571 => X"39",  -- 57
        2572 => X"39",  -- 57
        2573 => X"3A",  -- 58
        2574 => X"3C",  -- 60
        2575 => X"3D",  -- 61
        2576 => X"3D",  -- 61
        2577 => X"3D",  -- 61
        2578 => X"3D",  -- 61
        2579 => X"3D",  -- 61
        2580 => X"3D",  -- 61
        2581 => X"3D",  -- 61
        2582 => X"3D",  -- 61
        2583 => X"3D",  -- 61
        2584 => X"3C",  -- 60
        2585 => X"3D",  -- 61
        2586 => X"3E",  -- 62
        2587 => X"3E",  -- 62
        2588 => X"3E",  -- 62
        2589 => X"3E",  -- 62
        2590 => X"3E",  -- 62
        2591 => X"3E",  -- 62
        2592 => X"3D",  -- 61
        2593 => X"3C",  -- 60
        2594 => X"3B",  -- 59
        2595 => X"3A",  -- 58
        2596 => X"39",  -- 57
        2597 => X"38",  -- 56
        2598 => X"37",  -- 55
        2599 => X"37",  -- 55
        2600 => X"36",  -- 54
        2601 => X"36",  -- 54
        2602 => X"34",  -- 52
        2603 => X"33",  -- 51
        2604 => X"32",  -- 50
        2605 => X"31",  -- 49
        2606 => X"30",  -- 48
        2607 => X"30",  -- 48
        2608 => X"2E",  -- 46
        2609 => X"2E",  -- 46
        2610 => X"2E",  -- 46
        2611 => X"2E",  -- 46
        2612 => X"2C",  -- 44
        2613 => X"2B",  -- 43
        2614 => X"2A",  -- 42
        2615 => X"29",  -- 41
        2616 => X"28",  -- 40
        2617 => X"27",  -- 39
        2618 => X"25",  -- 37
        2619 => X"24",  -- 36
        2620 => X"24",  -- 36
        2621 => X"25",  -- 37
        2622 => X"25",  -- 37
        2623 => X"26",  -- 38
        2624 => X"29",  -- 41
        2625 => X"2C",  -- 44
        2626 => X"2E",  -- 46
        2627 => X"30",  -- 48
        2628 => X"31",  -- 49
        2629 => X"33",  -- 51
        2630 => X"37",  -- 55
        2631 => X"39",  -- 57
        2632 => X"3B",  -- 59
        2633 => X"3C",  -- 60
        2634 => X"3E",  -- 62
        2635 => X"41",  -- 65
        2636 => X"43",  -- 67
        2637 => X"45",  -- 69
        2638 => X"46",  -- 70
        2639 => X"46",  -- 70
        2640 => X"45",  -- 69
        2641 => X"43",  -- 67
        2642 => X"44",  -- 68
        2643 => X"48",  -- 72
        2644 => X"49",  -- 73
        2645 => X"44",  -- 68
        2646 => X"43",  -- 67
        2647 => X"46",  -- 70
        2648 => X"41",  -- 65
        2649 => X"66",  -- 102
        2650 => X"7B",  -- 123
        2651 => X"72",  -- 114
        2652 => X"67",  -- 103
        2653 => X"66",  -- 102
        2654 => X"5A",  -- 90
        2655 => X"43",  -- 67
        2656 => X"46",  -- 70
        2657 => X"4C",  -- 76
        2658 => X"68",  -- 104
        2659 => X"70",  -- 112
        2660 => X"5B",  -- 91
        2661 => X"60",  -- 96
        2662 => X"70",  -- 112
        2663 => X"68",  -- 104
        2664 => X"87",  -- 135
        2665 => X"7D",  -- 125
        2666 => X"76",  -- 118
        2667 => X"90",  -- 144
        2668 => X"8A",  -- 138
        2669 => X"8E",  -- 142
        2670 => X"7A",  -- 122
        2671 => X"70",  -- 112
        2672 => X"53",  -- 83
        2673 => X"44",  -- 68
        2674 => X"3B",  -- 59
        2675 => X"4D",  -- 77
        2676 => X"51",  -- 81
        2677 => X"3E",  -- 62
        2678 => X"40",  -- 64
        2679 => X"46",  -- 70
        2680 => X"56",  -- 86
        2681 => X"56",  -- 86
        2682 => X"46",  -- 70
        2683 => X"74",  -- 116
        2684 => X"85",  -- 133
        2685 => X"8E",  -- 142
        2686 => X"92",  -- 146
        2687 => X"8C",  -- 140
        2688 => X"98",  -- 152
        2689 => X"9C",  -- 156
        2690 => X"9A",  -- 154
        2691 => X"98",  -- 152
        2692 => X"9A",  -- 154
        2693 => X"9F",  -- 159
        2694 => X"99",  -- 153
        2695 => X"8E",  -- 142
        2696 => X"9A",  -- 154
        2697 => X"9E",  -- 158
        2698 => X"93",  -- 147
        2699 => X"8D",  -- 141
        2700 => X"96",  -- 150
        2701 => X"95",  -- 149
        2702 => X"8B",  -- 139
        2703 => X"8D",  -- 141
        2704 => X"A1",  -- 161
        2705 => X"8F",  -- 143
        2706 => X"8D",  -- 141
        2707 => X"9B",  -- 155
        2708 => X"9E",  -- 158
        2709 => X"90",  -- 144
        2710 => X"8B",  -- 139
        2711 => X"94",  -- 148
        2712 => X"A4",  -- 164
        2713 => X"9B",  -- 155
        2714 => X"9A",  -- 154
        2715 => X"A6",  -- 166
        2716 => X"A9",  -- 169
        2717 => X"A4",  -- 164
        2718 => X"A5",  -- 165
        2719 => X"AC",  -- 172
        2720 => X"B2",  -- 178
        2721 => X"AD",  -- 173
        2722 => X"A9",  -- 169
        2723 => X"A4",  -- 164
        2724 => X"9A",  -- 154
        2725 => X"89",  -- 137
        2726 => X"73",  -- 115
        2727 => X"65",  -- 101
        2728 => X"69",  -- 105
        2729 => X"6D",  -- 109
        2730 => X"6F",  -- 111
        2731 => X"6E",  -- 110
        2732 => X"6E",  -- 110
        2733 => X"75",  -- 117
        2734 => X"78",  -- 120
        2735 => X"75",  -- 117
        2736 => X"7E",  -- 126
        2737 => X"78",  -- 120
        2738 => X"7A",  -- 122
        2739 => X"83",  -- 131
        2740 => X"8B",  -- 139
        2741 => X"89",  -- 137
        2742 => X"84",  -- 132
        2743 => X"82",  -- 130
        2744 => X"89",  -- 137
        2745 => X"90",  -- 144
        2746 => X"8B",  -- 139
        2747 => X"8A",  -- 138
        2748 => X"94",  -- 148
        2749 => X"90",  -- 144
        2750 => X"86",  -- 134
        2751 => X"8B",  -- 139
        2752 => X"8F",  -- 143
        2753 => X"90",  -- 144
        2754 => X"93",  -- 147
        2755 => X"98",  -- 152
        2756 => X"9E",  -- 158
        2757 => X"A0",  -- 160
        2758 => X"9E",  -- 158
        2759 => X"9C",  -- 156
        2760 => X"A5",  -- 165
        2761 => X"A4",  -- 164
        2762 => X"A3",  -- 163
        2763 => X"A2",  -- 162
        2764 => X"A2",  -- 162
        2765 => X"A4",  -- 164
        2766 => X"A6",  -- 166
        2767 => X"A7",  -- 167
        2768 => X"A5",  -- 165
        2769 => X"AC",  -- 172
        2770 => X"B3",  -- 179
        2771 => X"B5",  -- 181
        2772 => X"B3",  -- 179
        2773 => X"B4",  -- 180
        2774 => X"B6",  -- 182
        2775 => X"B9",  -- 185
        2776 => X"B5",  -- 181
        2777 => X"B6",  -- 182
        2778 => X"B5",  -- 181
        2779 => X"AF",  -- 175
        2780 => X"AC",  -- 172
        2781 => X"AA",  -- 170
        2782 => X"A5",  -- 165
        2783 => X"9E",  -- 158
        2784 => X"95",  -- 149
        2785 => X"94",  -- 148
        2786 => X"95",  -- 149
        2787 => X"99",  -- 153
        2788 => X"98",  -- 152
        2789 => X"96",  -- 150
        2790 => X"98",  -- 152
        2791 => X"9C",  -- 156
        2792 => X"9B",  -- 155
        2793 => X"9E",  -- 158
        2794 => X"A1",  -- 161
        2795 => X"A0",  -- 160
        2796 => X"9D",  -- 157
        2797 => X"9B",  -- 155
        2798 => X"9E",  -- 158
        2799 => X"A2",  -- 162
        2800 => X"A5",  -- 165
        2801 => X"A3",  -- 163
        2802 => X"A3",  -- 163
        2803 => X"A4",  -- 164
        2804 => X"A8",  -- 168
        2805 => X"AC",  -- 172
        2806 => X"AE",  -- 174
        2807 => X"AE",  -- 174
        2808 => X"AD",  -- 173
        2809 => X"B3",  -- 179
        2810 => X"B4",  -- 180
        2811 => X"B1",  -- 177
        2812 => X"B1",  -- 177
        2813 => X"B5",  -- 181
        2814 => X"B5",  -- 181
        2815 => X"AE",  -- 174
        2816 => X"A9",  -- 169
        2817 => X"A2",  -- 162
        2818 => X"99",  -- 153
        2819 => X"95",  -- 149
        2820 => X"94",  -- 148
        2821 => X"94",  -- 148
        2822 => X"94",  -- 148
        2823 => X"92",  -- 146
        2824 => X"94",  -- 148
        2825 => X"98",  -- 152
        2826 => X"96",  -- 150
        2827 => X"8E",  -- 142
        2828 => X"85",  -- 133
        2829 => X"79",  -- 121
        2830 => X"6F",  -- 111
        2831 => X"65",  -- 101
        2832 => X"6A",  -- 106
        2833 => X"57",  -- 87
        2834 => X"4E",  -- 78
        2835 => X"4D",  -- 77
        2836 => X"46",  -- 70
        2837 => X"47",  -- 71
        2838 => X"50",  -- 80
        2839 => X"56",  -- 86
        2840 => X"55",  -- 85
        2841 => X"4E",  -- 78
        2842 => X"56",  -- 86
        2843 => X"6E",  -- 110
        2844 => X"7F",  -- 127
        2845 => X"88",  -- 136
        2846 => X"94",  -- 148
        2847 => X"A5",  -- 165
        2848 => X"AA",  -- 170
        2849 => X"AC",  -- 172
        2850 => X"B2",  -- 178
        2851 => X"BC",  -- 188
        2852 => X"BB",  -- 187
        2853 => X"B5",  -- 181
        2854 => X"B4",  -- 180
        2855 => X"B9",  -- 185
        2856 => X"B8",  -- 184
        2857 => X"B9",  -- 185
        2858 => X"BA",  -- 186
        2859 => X"BA",  -- 186
        2860 => X"BA",  -- 186
        2861 => X"B9",  -- 185
        2862 => X"BB",  -- 187
        2863 => X"BB",  -- 187
        2864 => X"B2",  -- 178
        2865 => X"B6",  -- 182
        2866 => X"B9",  -- 185
        2867 => X"B7",  -- 183
        2868 => X"B5",  -- 181
        2869 => X"B5",  -- 181
        2870 => X"B3",  -- 179
        2871 => X"AD",  -- 173
        2872 => X"B2",  -- 178
        2873 => X"AB",  -- 171
        2874 => X"A6",  -- 166
        2875 => X"A7",  -- 167
        2876 => X"AB",  -- 171
        2877 => X"AE",  -- 174
        2878 => X"B1",  -- 177
        2879 => X"B5",  -- 181
        2880 => X"3E",  -- 62
        2881 => X"3D",  -- 61
        2882 => X"3B",  -- 59
        2883 => X"3A",  -- 58
        2884 => X"38",  -- 56
        2885 => X"38",  -- 56
        2886 => X"39",  -- 57
        2887 => X"39",  -- 57
        2888 => X"39",  -- 57
        2889 => X"39",  -- 57
        2890 => X"39",  -- 57
        2891 => X"39",  -- 57
        2892 => X"3A",  -- 58
        2893 => X"3B",  -- 59
        2894 => X"3C",  -- 60
        2895 => X"3D",  -- 61
        2896 => X"3D",  -- 61
        2897 => X"3D",  -- 61
        2898 => X"3D",  -- 61
        2899 => X"3D",  -- 61
        2900 => X"3D",  -- 61
        2901 => X"3D",  -- 61
        2902 => X"3D",  -- 61
        2903 => X"3D",  -- 61
        2904 => X"3C",  -- 60
        2905 => X"3D",  -- 61
        2906 => X"3E",  -- 62
        2907 => X"3E",  -- 62
        2908 => X"3F",  -- 63
        2909 => X"3E",  -- 62
        2910 => X"3E",  -- 62
        2911 => X"3E",  -- 62
        2912 => X"3D",  -- 61
        2913 => X"3C",  -- 60
        2914 => X"3B",  -- 59
        2915 => X"3A",  -- 58
        2916 => X"3A",  -- 58
        2917 => X"38",  -- 56
        2918 => X"37",  -- 55
        2919 => X"37",  -- 55
        2920 => X"36",  -- 54
        2921 => X"36",  -- 54
        2922 => X"34",  -- 52
        2923 => X"33",  -- 51
        2924 => X"32",  -- 50
        2925 => X"31",  -- 49
        2926 => X"30",  -- 48
        2927 => X"30",  -- 48
        2928 => X"2F",  -- 47
        2929 => X"2F",  -- 47
        2930 => X"2E",  -- 46
        2931 => X"2E",  -- 46
        2932 => X"2D",  -- 45
        2933 => X"2B",  -- 43
        2934 => X"2A",  -- 42
        2935 => X"29",  -- 41
        2936 => X"28",  -- 40
        2937 => X"27",  -- 39
        2938 => X"26",  -- 38
        2939 => X"25",  -- 37
        2940 => X"24",  -- 36
        2941 => X"25",  -- 37
        2942 => X"26",  -- 38
        2943 => X"26",  -- 38
        2944 => X"2A",  -- 42
        2945 => X"2C",  -- 44
        2946 => X"2E",  -- 46
        2947 => X"30",  -- 48
        2948 => X"32",  -- 50
        2949 => X"34",  -- 52
        2950 => X"37",  -- 55
        2951 => X"3A",  -- 58
        2952 => X"3B",  -- 59
        2953 => X"3D",  -- 61
        2954 => X"3F",  -- 63
        2955 => X"41",  -- 65
        2956 => X"43",  -- 67
        2957 => X"45",  -- 69
        2958 => X"46",  -- 70
        2959 => X"47",  -- 71
        2960 => X"47",  -- 71
        2961 => X"45",  -- 69
        2962 => X"44",  -- 68
        2963 => X"46",  -- 70
        2964 => X"45",  -- 69
        2965 => X"45",  -- 69
        2966 => X"49",  -- 73
        2967 => X"4F",  -- 79
        2968 => X"50",  -- 80
        2969 => X"71",  -- 113
        2970 => X"8A",  -- 138
        2971 => X"84",  -- 132
        2972 => X"7C",  -- 124
        2973 => X"7B",  -- 123
        2974 => X"75",  -- 117
        2975 => X"68",  -- 104
        2976 => X"66",  -- 102
        2977 => X"68",  -- 104
        2978 => X"79",  -- 121
        2979 => X"77",  -- 119
        2980 => X"61",  -- 97
        2981 => X"68",  -- 104
        2982 => X"7E",  -- 126
        2983 => X"7E",  -- 126
        2984 => X"8D",  -- 141
        2985 => X"83",  -- 131
        2986 => X"7B",  -- 123
        2987 => X"8D",  -- 141
        2988 => X"88",  -- 136
        2989 => X"8C",  -- 140
        2990 => X"78",  -- 120
        2991 => X"69",  -- 105
        2992 => X"44",  -- 68
        2993 => X"39",  -- 57
        2994 => X"3F",  -- 63
        2995 => X"4C",  -- 76
        2996 => X"4B",  -- 75
        2997 => X"3E",  -- 62
        2998 => X"3E",  -- 62
        2999 => X"4E",  -- 78
        3000 => X"65",  -- 101
        3001 => X"61",  -- 97
        3002 => X"68",  -- 104
        3003 => X"7C",  -- 124
        3004 => X"89",  -- 137
        3005 => X"95",  -- 149
        3006 => X"90",  -- 144
        3007 => X"94",  -- 148
        3008 => X"96",  -- 150
        3009 => X"96",  -- 150
        3010 => X"98",  -- 152
        3011 => X"9A",  -- 154
        3012 => X"9E",  -- 158
        3013 => X"A0",  -- 160
        3014 => X"9A",  -- 154
        3015 => X"91",  -- 145
        3016 => X"93",  -- 147
        3017 => X"93",  -- 147
        3018 => X"93",  -- 147
        3019 => X"96",  -- 150
        3020 => X"8F",  -- 143
        3021 => X"80",  -- 128
        3022 => X"80",  -- 128
        3023 => X"91",  -- 145
        3024 => X"88",  -- 136
        3025 => X"8C",  -- 140
        3026 => X"91",  -- 145
        3027 => X"8E",  -- 142
        3028 => X"85",  -- 133
        3029 => X"82",  -- 130
        3030 => X"8C",  -- 140
        3031 => X"9A",  -- 154
        3032 => X"9A",  -- 154
        3033 => X"98",  -- 152
        3034 => X"9C",  -- 156
        3035 => X"A3",  -- 163
        3036 => X"A5",  -- 165
        3037 => X"A3",  -- 163
        3038 => X"A9",  -- 169
        3039 => X"B2",  -- 178
        3040 => X"B1",  -- 177
        3041 => X"AA",  -- 170
        3042 => X"A2",  -- 162
        3043 => X"9B",  -- 155
        3044 => X"94",  -- 148
        3045 => X"8A",  -- 138
        3046 => X"7E",  -- 126
        3047 => X"76",  -- 118
        3048 => X"64",  -- 100
        3049 => X"6A",  -- 106
        3050 => X"6E",  -- 110
        3051 => X"6D",  -- 109
        3052 => X"6E",  -- 110
        3053 => X"74",  -- 116
        3054 => X"7A",  -- 122
        3055 => X"7B",  -- 123
        3056 => X"80",  -- 128
        3057 => X"78",  -- 120
        3058 => X"75",  -- 117
        3059 => X"7A",  -- 122
        3060 => X"81",  -- 129
        3061 => X"83",  -- 131
        3062 => X"84",  -- 132
        3063 => X"86",  -- 134
        3064 => X"8B",  -- 139
        3065 => X"8D",  -- 141
        3066 => X"89",  -- 137
        3067 => X"88",  -- 136
        3068 => X"8F",  -- 143
        3069 => X"8F",  -- 143
        3070 => X"8C",  -- 140
        3071 => X"8F",  -- 143
        3072 => X"91",  -- 145
        3073 => X"91",  -- 145
        3074 => X"92",  -- 146
        3075 => X"96",  -- 150
        3076 => X"9B",  -- 155
        3077 => X"9C",  -- 156
        3078 => X"99",  -- 153
        3079 => X"97",  -- 151
        3080 => X"A3",  -- 163
        3081 => X"A3",  -- 163
        3082 => X"A2",  -- 162
        3083 => X"A1",  -- 161
        3084 => X"A1",  -- 161
        3085 => X"A2",  -- 162
        3086 => X"A3",  -- 163
        3087 => X"A4",  -- 164
        3088 => X"A7",  -- 167
        3089 => X"AA",  -- 170
        3090 => X"AE",  -- 174
        3091 => X"B2",  -- 178
        3092 => X"B3",  -- 179
        3093 => X"B6",  -- 182
        3094 => X"B6",  -- 182
        3095 => X"B7",  -- 183
        3096 => X"B7",  -- 183
        3097 => X"B7",  -- 183
        3098 => X"B4",  -- 180
        3099 => X"AE",  -- 174
        3100 => X"AD",  -- 173
        3101 => X"AB",  -- 171
        3102 => X"A5",  -- 165
        3103 => X"9D",  -- 157
        3104 => X"99",  -- 153
        3105 => X"95",  -- 149
        3106 => X"94",  -- 148
        3107 => X"93",  -- 147
        3108 => X"90",  -- 144
        3109 => X"8D",  -- 141
        3110 => X"90",  -- 144
        3111 => X"94",  -- 148
        3112 => X"9B",  -- 155
        3113 => X"9C",  -- 156
        3114 => X"9F",  -- 159
        3115 => X"A0",  -- 160
        3116 => X"A2",  -- 162
        3117 => X"A3",  -- 163
        3118 => X"A4",  -- 164
        3119 => X"A5",  -- 165
        3120 => X"A8",  -- 168
        3121 => X"A8",  -- 168
        3122 => X"A7",  -- 167
        3123 => X"A5",  -- 165
        3124 => X"A4",  -- 164
        3125 => X"A5",  -- 165
        3126 => X"AA",  -- 170
        3127 => X"AC",  -- 172
        3128 => X"B0",  -- 176
        3129 => X"B2",  -- 178
        3130 => X"B2",  -- 178
        3131 => X"B1",  -- 177
        3132 => X"B2",  -- 178
        3133 => X"B5",  -- 181
        3134 => X"B7",  -- 183
        3135 => X"B6",  -- 182
        3136 => X"AF",  -- 175
        3137 => X"A7",  -- 167
        3138 => X"9B",  -- 155
        3139 => X"96",  -- 150
        3140 => X"94",  -- 148
        3141 => X"95",  -- 149
        3142 => X"96",  -- 150
        3143 => X"95",  -- 149
        3144 => X"98",  -- 152
        3145 => X"96",  -- 150
        3146 => X"93",  -- 147
        3147 => X"8F",  -- 143
        3148 => X"8B",  -- 139
        3149 => X"83",  -- 131
        3150 => X"75",  -- 117
        3151 => X"68",  -- 104
        3152 => X"60",  -- 96
        3153 => X"58",  -- 88
        3154 => X"59",  -- 89
        3155 => X"59",  -- 89
        3156 => X"51",  -- 81
        3157 => X"4F",  -- 79
        3158 => X"55",  -- 85
        3159 => X"56",  -- 86
        3160 => X"46",  -- 70
        3161 => X"42",  -- 66
        3162 => X"4C",  -- 76
        3163 => X"61",  -- 97
        3164 => X"72",  -- 114
        3165 => X"79",  -- 121
        3166 => X"84",  -- 132
        3167 => X"93",  -- 147
        3168 => X"9E",  -- 158
        3169 => X"A6",  -- 166
        3170 => X"B4",  -- 180
        3171 => X"BB",  -- 187
        3172 => X"B9",  -- 185
        3173 => X"B5",  -- 181
        3174 => X"B5",  -- 181
        3175 => X"B8",  -- 184
        3176 => X"BA",  -- 186
        3177 => X"B9",  -- 185
        3178 => X"B6",  -- 182
        3179 => X"B3",  -- 179
        3180 => X"B3",  -- 179
        3181 => X"B4",  -- 180
        3182 => X"B8",  -- 184
        3183 => X"BC",  -- 188
        3184 => X"B7",  -- 183
        3185 => X"BB",  -- 187
        3186 => X"BC",  -- 188
        3187 => X"B8",  -- 184
        3188 => X"B6",  -- 182
        3189 => X"B8",  -- 184
        3190 => X"B7",  -- 183
        3191 => X"B3",  -- 179
        3192 => X"AC",  -- 172
        3193 => X"A8",  -- 168
        3194 => X"A7",  -- 167
        3195 => X"AB",  -- 171
        3196 => X"AE",  -- 174
        3197 => X"AE",  -- 174
        3198 => X"B1",  -- 177
        3199 => X"B4",  -- 180
        3200 => X"3F",  -- 63
        3201 => X"3E",  -- 62
        3202 => X"3D",  -- 61
        3203 => X"3B",  -- 59
        3204 => X"39",  -- 57
        3205 => X"39",  -- 57
        3206 => X"3A",  -- 58
        3207 => X"3A",  -- 58
        3208 => X"3A",  -- 58
        3209 => X"39",  -- 57
        3210 => X"39",  -- 57
        3211 => X"39",  -- 57
        3212 => X"3A",  -- 58
        3213 => X"3B",  -- 59
        3214 => X"3D",  -- 61
        3215 => X"3D",  -- 61
        3216 => X"3D",  -- 61
        3217 => X"3D",  -- 61
        3218 => X"3D",  -- 61
        3219 => X"3D",  -- 61
        3220 => X"3D",  -- 61
        3221 => X"3D",  -- 61
        3222 => X"3D",  -- 61
        3223 => X"3D",  -- 61
        3224 => X"3D",  -- 61
        3225 => X"3D",  -- 61
        3226 => X"3E",  -- 62
        3227 => X"3F",  -- 63
        3228 => X"3F",  -- 63
        3229 => X"3F",  -- 63
        3230 => X"3E",  -- 62
        3231 => X"3E",  -- 62
        3232 => X"3D",  -- 61
        3233 => X"3C",  -- 60
        3234 => X"3B",  -- 59
        3235 => X"3A",  -- 58
        3236 => X"3A",  -- 58
        3237 => X"39",  -- 57
        3238 => X"38",  -- 56
        3239 => X"37",  -- 55
        3240 => X"37",  -- 55
        3241 => X"36",  -- 54
        3242 => X"34",  -- 52
        3243 => X"33",  -- 51
        3244 => X"32",  -- 50
        3245 => X"31",  -- 49
        3246 => X"30",  -- 48
        3247 => X"30",  -- 48
        3248 => X"2F",  -- 47
        3249 => X"2F",  -- 47
        3250 => X"2F",  -- 47
        3251 => X"2E",  -- 46
        3252 => X"2D",  -- 45
        3253 => X"2B",  -- 43
        3254 => X"2A",  -- 42
        3255 => X"29",  -- 41
        3256 => X"28",  -- 40
        3257 => X"27",  -- 39
        3258 => X"26",  -- 38
        3259 => X"25",  -- 37
        3260 => X"25",  -- 37
        3261 => X"25",  -- 37
        3262 => X"26",  -- 38
        3263 => X"27",  -- 39
        3264 => X"2A",  -- 42
        3265 => X"2C",  -- 44
        3266 => X"2F",  -- 47
        3267 => X"31",  -- 49
        3268 => X"32",  -- 50
        3269 => X"34",  -- 52
        3270 => X"38",  -- 56
        3271 => X"3A",  -- 58
        3272 => X"3C",  -- 60
        3273 => X"3D",  -- 61
        3274 => X"3F",  -- 63
        3275 => X"42",  -- 66
        3276 => X"44",  -- 68
        3277 => X"46",  -- 70
        3278 => X"47",  -- 71
        3279 => X"48",  -- 72
        3280 => X"47",  -- 71
        3281 => X"47",  -- 71
        3282 => X"48",  -- 72
        3283 => X"47",  -- 71
        3284 => X"48",  -- 72
        3285 => X"4A",  -- 74
        3286 => X"53",  -- 83
        3287 => X"5D",  -- 93
        3288 => X"66",  -- 102
        3289 => X"81",  -- 129
        3290 => X"95",  -- 149
        3291 => X"95",  -- 149
        3292 => X"8D",  -- 141
        3293 => X"8D",  -- 141
        3294 => X"8C",  -- 140
        3295 => X"8A",  -- 138
        3296 => X"87",  -- 135
        3297 => X"86",  -- 134
        3298 => X"8F",  -- 143
        3299 => X"86",  -- 134
        3300 => X"70",  -- 112
        3301 => X"75",  -- 117
        3302 => X"8D",  -- 141
        3303 => X"91",  -- 145
        3304 => X"91",  -- 145
        3305 => X"87",  -- 135
        3306 => X"7F",  -- 127
        3307 => X"87",  -- 135
        3308 => X"81",  -- 129
        3309 => X"84",  -- 132
        3310 => X"70",  -- 112
        3311 => X"5B",  -- 91
        3312 => X"38",  -- 56
        3313 => X"31",  -- 49
        3314 => X"48",  -- 72
        3315 => X"4A",  -- 74
        3316 => X"44",  -- 68
        3317 => X"40",  -- 64
        3318 => X"43",  -- 67
        3319 => X"65",  -- 101
        3320 => X"77",  -- 119
        3321 => X"72",  -- 114
        3322 => X"8D",  -- 141
        3323 => X"86",  -- 134
        3324 => X"8F",  -- 143
        3325 => X"98",  -- 152
        3326 => X"8E",  -- 142
        3327 => X"98",  -- 152
        3328 => X"97",  -- 151
        3329 => X"94",  -- 148
        3330 => X"94",  -- 148
        3331 => X"9C",  -- 156
        3332 => X"A0",  -- 160
        3333 => X"9B",  -- 155
        3334 => X"96",  -- 150
        3335 => X"92",  -- 146
        3336 => X"8E",  -- 142
        3337 => X"8A",  -- 138
        3338 => X"8D",  -- 141
        3339 => X"8D",  -- 141
        3340 => X"80",  -- 128
        3341 => X"79",  -- 121
        3342 => X"83",  -- 131
        3343 => X"8D",  -- 141
        3344 => X"77",  -- 119
        3345 => X"85",  -- 133
        3346 => X"8B",  -- 139
        3347 => X"7D",  -- 125
        3348 => X"73",  -- 115
        3349 => X"79",  -- 121
        3350 => X"89",  -- 137
        3351 => X"92",  -- 146
        3352 => X"93",  -- 147
        3353 => X"99",  -- 153
        3354 => X"9F",  -- 159
        3355 => X"9F",  -- 159
        3356 => X"9C",  -- 156
        3357 => X"9E",  -- 158
        3358 => X"A5",  -- 165
        3359 => X"AC",  -- 172
        3360 => X"A4",  -- 164
        3361 => X"A5",  -- 165
        3362 => X"A7",  -- 167
        3363 => X"A4",  -- 164
        3364 => X"9A",  -- 154
        3365 => X"8B",  -- 139
        3366 => X"79",  -- 121
        3367 => X"6C",  -- 108
        3368 => X"64",  -- 100
        3369 => X"68",  -- 104
        3370 => X"6C",  -- 108
        3371 => X"6B",  -- 107
        3372 => X"6D",  -- 109
        3373 => X"73",  -- 115
        3374 => X"78",  -- 120
        3375 => X"7A",  -- 122
        3376 => X"77",  -- 119
        3377 => X"72",  -- 114
        3378 => X"71",  -- 113
        3379 => X"75",  -- 117
        3380 => X"7D",  -- 125
        3381 => X"80",  -- 128
        3382 => X"83",  -- 131
        3383 => X"86",  -- 134
        3384 => X"8B",  -- 139
        3385 => X"85",  -- 133
        3386 => X"86",  -- 134
        3387 => X"88",  -- 136
        3388 => X"87",  -- 135
        3389 => X"8B",  -- 139
        3390 => X"90",  -- 144
        3391 => X"8F",  -- 143
        3392 => X"8B",  -- 139
        3393 => X"8B",  -- 139
        3394 => X"8E",  -- 142
        3395 => X"93",  -- 147
        3396 => X"97",  -- 151
        3397 => X"9A",  -- 154
        3398 => X"9C",  -- 156
        3399 => X"9C",  -- 156
        3400 => X"A1",  -- 161
        3401 => X"A1",  -- 161
        3402 => X"A2",  -- 162
        3403 => X"A2",  -- 162
        3404 => X"A1",  -- 161
        3405 => X"A1",  -- 161
        3406 => X"A2",  -- 162
        3407 => X"A4",  -- 164
        3408 => X"A9",  -- 169
        3409 => X"A9",  -- 169
        3410 => X"AA",  -- 170
        3411 => X"AF",  -- 175
        3412 => X"B3",  -- 179
        3413 => X"B7",  -- 183
        3414 => X"B6",  -- 182
        3415 => X"B5",  -- 181
        3416 => X"B9",  -- 185
        3417 => X"B7",  -- 183
        3418 => X"B4",  -- 180
        3419 => X"AE",  -- 174
        3420 => X"AE",  -- 174
        3421 => X"AC",  -- 172
        3422 => X"A6",  -- 166
        3423 => X"9C",  -- 156
        3424 => X"9B",  -- 155
        3425 => X"96",  -- 150
        3426 => X"93",  -- 147
        3427 => X"92",  -- 146
        3428 => X"91",  -- 145
        3429 => X"90",  -- 144
        3430 => X"95",  -- 149
        3431 => X"9A",  -- 154
        3432 => X"9A",  -- 154
        3433 => X"9A",  -- 154
        3434 => X"9B",  -- 155
        3435 => X"A0",  -- 160
        3436 => X"A5",  -- 165
        3437 => X"A8",  -- 168
        3438 => X"A8",  -- 168
        3439 => X"A6",  -- 166
        3440 => X"A6",  -- 166
        3441 => X"A8",  -- 168
        3442 => X"A9",  -- 169
        3443 => X"A5",  -- 165
        3444 => X"A1",  -- 161
        3445 => X"A1",  -- 161
        3446 => X"A6",  -- 166
        3447 => X"AC",  -- 172
        3448 => X"B0",  -- 176
        3449 => X"AD",  -- 173
        3450 => X"AE",  -- 174
        3451 => X"B0",  -- 176
        3452 => X"B1",  -- 177
        3453 => X"B3",  -- 179
        3454 => X"B7",  -- 183
        3455 => X"BC",  -- 188
        3456 => X"B5",  -- 181
        3457 => X"AD",  -- 173
        3458 => X"A1",  -- 161
        3459 => X"9A",  -- 154
        3460 => X"98",  -- 152
        3461 => X"98",  -- 152
        3462 => X"99",  -- 153
        3463 => X"9A",  -- 154
        3464 => X"9A",  -- 154
        3465 => X"95",  -- 149
        3466 => X"90",  -- 144
        3467 => X"8F",  -- 143
        3468 => X"91",  -- 145
        3469 => X"8D",  -- 141
        3470 => X"7D",  -- 125
        3471 => X"6D",  -- 109
        3472 => X"67",  -- 103
        3473 => X"66",  -- 102
        3474 => X"6A",  -- 106
        3475 => X"62",  -- 98
        3476 => X"55",  -- 85
        3477 => X"55",  -- 85
        3478 => X"58",  -- 88
        3479 => X"51",  -- 81
        3480 => X"42",  -- 66
        3481 => X"45",  -- 69
        3482 => X"52",  -- 82
        3483 => X"66",  -- 102
        3484 => X"6D",  -- 109
        3485 => X"6D",  -- 109
        3486 => X"71",  -- 113
        3487 => X"7B",  -- 123
        3488 => X"86",  -- 134
        3489 => X"98",  -- 152
        3490 => X"AC",  -- 172
        3491 => X"B5",  -- 181
        3492 => X"B6",  -- 182
        3493 => X"B8",  -- 184
        3494 => X"BB",  -- 187
        3495 => X"BC",  -- 188
        3496 => X"B7",  -- 183
        3497 => X"B6",  -- 182
        3498 => X"B6",  -- 182
        3499 => X"B5",  -- 181
        3500 => X"B4",  -- 180
        3501 => X"B6",  -- 182
        3502 => X"B8",  -- 184
        3503 => X"BC",  -- 188
        3504 => X"BC",  -- 188
        3505 => X"BC",  -- 188
        3506 => X"BA",  -- 186
        3507 => X"B6",  -- 182
        3508 => X"B5",  -- 181
        3509 => X"B7",  -- 183
        3510 => X"B7",  -- 183
        3511 => X"B6",  -- 182
        3512 => X"AC",  -- 172
        3513 => X"AB",  -- 171
        3514 => X"AD",  -- 173
        3515 => X"B1",  -- 177
        3516 => X"B1",  -- 177
        3517 => X"AE",  -- 174
        3518 => X"AF",  -- 175
        3519 => X"B3",  -- 179
        3520 => X"41",  -- 65
        3521 => X"40",  -- 64
        3522 => X"3E",  -- 62
        3523 => X"3C",  -- 60
        3524 => X"3A",  -- 58
        3525 => X"3A",  -- 58
        3526 => X"3B",  -- 59
        3527 => X"3B",  -- 59
        3528 => X"3A",  -- 58
        3529 => X"3A",  -- 58
        3530 => X"3A",  -- 58
        3531 => X"3A",  -- 58
        3532 => X"3A",  -- 58
        3533 => X"3B",  -- 59
        3534 => X"3D",  -- 61
        3535 => X"3E",  -- 62
        3536 => X"3E",  -- 62
        3537 => X"3E",  -- 62
        3538 => X"3E",  -- 62
        3539 => X"3E",  -- 62
        3540 => X"3E",  -- 62
        3541 => X"3E",  -- 62
        3542 => X"3E",  -- 62
        3543 => X"3E",  -- 62
        3544 => X"3D",  -- 61
        3545 => X"3D",  -- 61
        3546 => X"3E",  -- 62
        3547 => X"3F",  -- 63
        3548 => X"3F",  -- 63
        3549 => X"3F",  -- 63
        3550 => X"3F",  -- 63
        3551 => X"3E",  -- 62
        3552 => X"3D",  -- 61
        3553 => X"3D",  -- 61
        3554 => X"3C",  -- 60
        3555 => X"3B",  -- 59
        3556 => X"3A",  -- 58
        3557 => X"39",  -- 57
        3558 => X"38",  -- 56
        3559 => X"37",  -- 55
        3560 => X"37",  -- 55
        3561 => X"36",  -- 54
        3562 => X"35",  -- 53
        3563 => X"34",  -- 52
        3564 => X"33",  -- 51
        3565 => X"31",  -- 49
        3566 => X"31",  -- 49
        3567 => X"30",  -- 48
        3568 => X"2F",  -- 47
        3569 => X"2F",  -- 47
        3570 => X"2F",  -- 47
        3571 => X"2E",  -- 46
        3572 => X"2D",  -- 45
        3573 => X"2C",  -- 44
        3574 => X"2A",  -- 42
        3575 => X"2A",  -- 42
        3576 => X"29",  -- 41
        3577 => X"28",  -- 40
        3578 => X"27",  -- 39
        3579 => X"26",  -- 38
        3580 => X"25",  -- 37
        3581 => X"26",  -- 38
        3582 => X"27",  -- 39
        3583 => X"28",  -- 40
        3584 => X"2A",  -- 42
        3585 => X"2C",  -- 44
        3586 => X"2F",  -- 47
        3587 => X"31",  -- 49
        3588 => X"33",  -- 51
        3589 => X"35",  -- 53
        3590 => X"39",  -- 57
        3591 => X"3B",  -- 59
        3592 => X"3D",  -- 61
        3593 => X"3E",  -- 62
        3594 => X"40",  -- 64
        3595 => X"43",  -- 67
        3596 => X"45",  -- 69
        3597 => X"47",  -- 71
        3598 => X"48",  -- 72
        3599 => X"49",  -- 73
        3600 => X"45",  -- 69
        3601 => X"49",  -- 73
        3602 => X"4B",  -- 75
        3603 => X"4C",  -- 76
        3604 => X"4F",  -- 79
        3605 => X"58",  -- 88
        3606 => X"65",  -- 101
        3607 => X"72",  -- 114
        3608 => X"85",  -- 133
        3609 => X"91",  -- 145
        3610 => X"9B",  -- 155
        3611 => X"9E",  -- 158
        3612 => X"9A",  -- 154
        3613 => X"96",  -- 150
        3614 => X"96",  -- 150
        3615 => X"99",  -- 153
        3616 => X"92",  -- 146
        3617 => X"95",  -- 149
        3618 => X"9B",  -- 155
        3619 => X"95",  -- 149
        3620 => X"85",  -- 133
        3621 => X"87",  -- 135
        3622 => X"93",  -- 147
        3623 => X"92",  -- 146
        3624 => X"90",  -- 144
        3625 => X"88",  -- 136
        3626 => X"83",  -- 131
        3627 => X"80",  -- 128
        3628 => X"7A",  -- 122
        3629 => X"78",  -- 120
        3630 => X"64",  -- 100
        3631 => X"49",  -- 73
        3632 => X"33",  -- 51
        3633 => X"32",  -- 50
        3634 => X"56",  -- 86
        3635 => X"51",  -- 81
        3636 => X"47",  -- 71
        3637 => X"4E",  -- 78
        3638 => X"51",  -- 81
        3639 => X"7F",  -- 127
        3640 => X"7F",  -- 127
        3641 => X"82",  -- 130
        3642 => X"9A",  -- 154
        3643 => X"8C",  -- 140
        3644 => X"95",  -- 149
        3645 => X"93",  -- 147
        3646 => X"93",  -- 147
        3647 => X"94",  -- 148
        3648 => X"9C",  -- 156
        3649 => X"95",  -- 149
        3650 => X"92",  -- 146
        3651 => X"99",  -- 153
        3652 => X"99",  -- 153
        3653 => X"92",  -- 146
        3654 => X"8D",  -- 141
        3655 => X"8F",  -- 143
        3656 => X"8C",  -- 140
        3657 => X"84",  -- 132
        3658 => X"80",  -- 128
        3659 => X"71",  -- 113
        3660 => X"6D",  -- 109
        3661 => X"82",  -- 130
        3662 => X"8C",  -- 140
        3663 => X"78",  -- 120
        3664 => X"6D",  -- 109
        3665 => X"70",  -- 112
        3666 => X"6E",  -- 110
        3667 => X"69",  -- 105
        3668 => X"6F",  -- 111
        3669 => X"7D",  -- 125
        3670 => X"83",  -- 131
        3671 => X"81",  -- 129
        3672 => X"82",  -- 130
        3673 => X"8E",  -- 142
        3674 => X"97",  -- 151
        3675 => X"96",  -- 150
        3676 => X"96",  -- 150
        3677 => X"9C",  -- 156
        3678 => X"A1",  -- 161
        3679 => X"A0",  -- 160
        3680 => X"B0",  -- 176
        3681 => X"AB",  -- 171
        3682 => X"A0",  -- 160
        3683 => X"94",  -- 148
        3684 => X"8A",  -- 138
        3685 => X"81",  -- 129
        3686 => X"7B",  -- 123
        3687 => X"7A",  -- 122
        3688 => X"6C",  -- 108
        3689 => X"6B",  -- 107
        3690 => X"6A",  -- 106
        3691 => X"6B",  -- 107
        3692 => X"6E",  -- 110
        3693 => X"71",  -- 113
        3694 => X"72",  -- 114
        3695 => X"72",  -- 114
        3696 => X"69",  -- 105
        3697 => X"6B",  -- 107
        3698 => X"71",  -- 113
        3699 => X"79",  -- 121
        3700 => X"80",  -- 128
        3701 => X"82",  -- 130
        3702 => X"81",  -- 129
        3703 => X"81",  -- 129
        3704 => X"87",  -- 135
        3705 => X"7D",  -- 125
        3706 => X"82",  -- 130
        3707 => X"87",  -- 135
        3708 => X"82",  -- 130
        3709 => X"89",  -- 137
        3710 => X"91",  -- 145
        3711 => X"89",  -- 137
        3712 => X"87",  -- 135
        3713 => X"89",  -- 137
        3714 => X"8C",  -- 140
        3715 => X"90",  -- 144
        3716 => X"94",  -- 148
        3717 => X"99",  -- 153
        3718 => X"9B",  -- 155
        3719 => X"9D",  -- 157
        3720 => X"9D",  -- 157
        3721 => X"A0",  -- 160
        3722 => X"A2",  -- 162
        3723 => X"A3",  -- 163
        3724 => X"A3",  -- 163
        3725 => X"A3",  -- 163
        3726 => X"A5",  -- 165
        3727 => X"A7",  -- 167
        3728 => X"A9",  -- 169
        3729 => X"AA",  -- 170
        3730 => X"AC",  -- 172
        3731 => X"AF",  -- 175
        3732 => X"B2",  -- 178
        3733 => X"B6",  -- 182
        3734 => X"B7",  -- 183
        3735 => X"B7",  -- 183
        3736 => X"BB",  -- 187
        3737 => X"B8",  -- 184
        3738 => X"B4",  -- 180
        3739 => X"AE",  -- 174
        3740 => X"AF",  -- 175
        3741 => X"AE",  -- 174
        3742 => X"A6",  -- 166
        3743 => X"9C",  -- 156
        3744 => X"9B",  -- 155
        3745 => X"96",  -- 150
        3746 => X"94",  -- 148
        3747 => X"95",  -- 149
        3748 => X"94",  -- 148
        3749 => X"93",  -- 147
        3750 => X"98",  -- 152
        3751 => X"9E",  -- 158
        3752 => X"99",  -- 153
        3753 => X"9A",  -- 154
        3754 => X"9C",  -- 156
        3755 => X"9F",  -- 159
        3756 => X"A3",  -- 163
        3757 => X"A5",  -- 165
        3758 => X"A5",  -- 165
        3759 => X"A4",  -- 164
        3760 => X"A0",  -- 160
        3761 => X"A3",  -- 163
        3762 => X"A6",  -- 166
        3763 => X"A5",  -- 165
        3764 => X"A4",  -- 164
        3765 => X"A4",  -- 164
        3766 => X"A8",  -- 168
        3767 => X"AC",  -- 172
        3768 => X"AD",  -- 173
        3769 => X"A8",  -- 168
        3770 => X"A9",  -- 169
        3771 => X"B0",  -- 176
        3772 => X"B2",  -- 178
        3773 => X"B1",  -- 177
        3774 => X"B5",  -- 181
        3775 => X"BC",  -- 188
        3776 => X"B9",  -- 185
        3777 => X"B2",  -- 178
        3778 => X"AA",  -- 170
        3779 => X"A1",  -- 161
        3780 => X"9E",  -- 158
        3781 => X"9D",  -- 157
        3782 => X"9C",  -- 156
        3783 => X"9C",  -- 156
        3784 => X"9A",  -- 154
        3785 => X"97",  -- 151
        3786 => X"92",  -- 146
        3787 => X"91",  -- 145
        3788 => X"94",  -- 148
        3789 => X"92",  -- 146
        3790 => X"85",  -- 133
        3791 => X"76",  -- 118
        3792 => X"7D",  -- 125
        3793 => X"7B",  -- 123
        3794 => X"76",  -- 118
        3795 => X"67",  -- 103
        3796 => X"58",  -- 88
        3797 => X"5B",  -- 91
        3798 => X"5A",  -- 90
        3799 => X"4E",  -- 78
        3800 => X"44",  -- 68
        3801 => X"52",  -- 82
        3802 => X"66",  -- 102
        3803 => X"73",  -- 115
        3804 => X"6E",  -- 110
        3805 => X"63",  -- 99
        3806 => X"5F",  -- 95
        3807 => X"63",  -- 99
        3808 => X"73",  -- 115
        3809 => X"89",  -- 137
        3810 => X"9F",  -- 159
        3811 => X"AA",  -- 170
        3812 => X"B0",  -- 176
        3813 => X"B7",  -- 183
        3814 => X"BB",  -- 187
        3815 => X"B9",  -- 185
        3816 => X"B1",  -- 177
        3817 => X"B6",  -- 182
        3818 => X"BB",  -- 187
        3819 => X"BE",  -- 190
        3820 => X"BF",  -- 191
        3821 => X"BE",  -- 190
        3822 => X"BE",  -- 190
        3823 => X"BE",  -- 190
        3824 => X"BD",  -- 189
        3825 => X"BB",  -- 187
        3826 => X"B7",  -- 183
        3827 => X"B2",  -- 178
        3828 => X"B1",  -- 177
        3829 => X"B3",  -- 179
        3830 => X"B4",  -- 180
        3831 => X"B5",  -- 181
        3832 => X"B4",  -- 180
        3833 => X"B4",  -- 180
        3834 => X"B5",  -- 181
        3835 => X"B7",  -- 183
        3836 => X"B3",  -- 179
        3837 => X"AF",  -- 175
        3838 => X"AF",  -- 175
        3839 => X"B3",  -- 179
        3840 => X"42",  -- 66
        3841 => X"41",  -- 65
        3842 => X"3F",  -- 63
        3843 => X"3D",  -- 61
        3844 => X"3B",  -- 59
        3845 => X"3B",  -- 59
        3846 => X"3B",  -- 59
        3847 => X"3B",  -- 59
        3848 => X"3A",  -- 58
        3849 => X"3A",  -- 58
        3850 => X"3A",  -- 58
        3851 => X"3A",  -- 58
        3852 => X"3B",  -- 59
        3853 => X"3B",  -- 59
        3854 => X"3D",  -- 61
        3855 => X"3E",  -- 62
        3856 => X"3E",  -- 62
        3857 => X"3E",  -- 62
        3858 => X"3E",  -- 62
        3859 => X"3E",  -- 62
        3860 => X"3E",  -- 62
        3861 => X"3E",  -- 62
        3862 => X"3E",  -- 62
        3863 => X"3E",  -- 62
        3864 => X"3D",  -- 61
        3865 => X"3E",  -- 62
        3866 => X"3F",  -- 63
        3867 => X"3F",  -- 63
        3868 => X"3F",  -- 63
        3869 => X"3F",  -- 63
        3870 => X"3F",  -- 63
        3871 => X"3F",  -- 63
        3872 => X"3E",  -- 62
        3873 => X"3D",  -- 61
        3874 => X"3C",  -- 60
        3875 => X"3B",  -- 59
        3876 => X"3A",  -- 58
        3877 => X"39",  -- 57
        3878 => X"38",  -- 56
        3879 => X"38",  -- 56
        3880 => X"37",  -- 55
        3881 => X"37",  -- 55
        3882 => X"35",  -- 53
        3883 => X"34",  -- 52
        3884 => X"33",  -- 51
        3885 => X"32",  -- 50
        3886 => X"31",  -- 49
        3887 => X"31",  -- 49
        3888 => X"30",  -- 48
        3889 => X"30",  -- 48
        3890 => X"2F",  -- 47
        3891 => X"2F",  -- 47
        3892 => X"2E",  -- 46
        3893 => X"2C",  -- 44
        3894 => X"2B",  -- 43
        3895 => X"2A",  -- 42
        3896 => X"2A",  -- 42
        3897 => X"29",  -- 41
        3898 => X"27",  -- 39
        3899 => X"26",  -- 38
        3900 => X"26",  -- 38
        3901 => X"27",  -- 39
        3902 => X"28",  -- 40
        3903 => X"28",  -- 40
        3904 => X"2A",  -- 42
        3905 => X"2C",  -- 44
        3906 => X"2F",  -- 47
        3907 => X"32",  -- 50
        3908 => X"34",  -- 52
        3909 => X"36",  -- 54
        3910 => X"3A",  -- 58
        3911 => X"3D",  -- 61
        3912 => X"3E",  -- 62
        3913 => X"3F",  -- 63
        3914 => X"41",  -- 65
        3915 => X"44",  -- 68
        3916 => X"46",  -- 70
        3917 => X"48",  -- 72
        3918 => X"49",  -- 73
        3919 => X"4A",  -- 74
        3920 => X"48",  -- 72
        3921 => X"4B",  -- 75
        3922 => X"4A",  -- 74
        3923 => X"4B",  -- 75
        3924 => X"52",  -- 82
        3925 => X"64",  -- 100
        3926 => X"7B",  -- 123
        3927 => X"8D",  -- 141
        3928 => X"A1",  -- 161
        3929 => X"9F",  -- 159
        3930 => X"9E",  -- 158
        3931 => X"A2",  -- 162
        3932 => X"A2",  -- 162
        3933 => X"A0",  -- 160
        3934 => X"9D",  -- 157
        3935 => X"9C",  -- 156
        3936 => X"94",  -- 148
        3937 => X"96",  -- 150
        3938 => X"9C",  -- 156
        3939 => X"9B",  -- 155
        3940 => X"96",  -- 150
        3941 => X"95",  -- 149
        3942 => X"95",  -- 149
        3943 => X"8D",  -- 141
        3944 => X"8C",  -- 140
        3945 => X"86",  -- 134
        3946 => X"84",  -- 132
        3947 => X"7B",  -- 123
        3948 => X"73",  -- 115
        3949 => X"6B",  -- 107
        3950 => X"57",  -- 87
        3951 => X"3B",  -- 59
        3952 => X"31",  -- 49
        3953 => X"3A",  -- 58
        3954 => X"67",  -- 103
        3955 => X"65",  -- 101
        3956 => X"5B",  -- 91
        3957 => X"60",  -- 96
        3958 => X"61",  -- 97
        3959 => X"8B",  -- 139
        3960 => X"81",  -- 129
        3961 => X"8C",  -- 140
        3962 => X"92",  -- 146
        3963 => X"8F",  -- 143
        3964 => X"9A",  -- 154
        3965 => X"8C",  -- 140
        3966 => X"9A",  -- 154
        3967 => X"8F",  -- 143
        3968 => X"9C",  -- 156
        3969 => X"94",  -- 148
        3970 => X"8F",  -- 143
        3971 => X"91",  -- 145
        3972 => X"8F",  -- 143
        3973 => X"88",  -- 136
        3974 => X"85",  -- 133
        3975 => X"88",  -- 136
        3976 => X"81",  -- 129
        3977 => X"77",  -- 119
        3978 => X"6F",  -- 111
        3979 => X"65",  -- 101
        3980 => X"64",  -- 100
        3981 => X"7A",  -- 122
        3982 => X"7B",  -- 123
        3983 => X"5F",  -- 95
        3984 => X"5C",  -- 92
        3985 => X"53",  -- 83
        3986 => X"50",  -- 80
        3987 => X"5A",  -- 90
        3988 => X"6A",  -- 106
        3989 => X"73",  -- 115
        3990 => X"70",  -- 112
        3991 => X"6B",  -- 107
        3992 => X"67",  -- 103
        3993 => X"74",  -- 116
        3994 => X"82",  -- 130
        3995 => X"87",  -- 135
        3996 => X"8E",  -- 142
        3997 => X"99",  -- 153
        3998 => X"9F",  -- 159
        3999 => X"9C",  -- 156
        4000 => X"A8",  -- 168
        4001 => X"A6",  -- 166
        4002 => X"9F",  -- 159
        4003 => X"97",  -- 151
        4004 => X"8F",  -- 143
        4005 => X"85",  -- 133
        4006 => X"7F",  -- 127
        4007 => X"7C",  -- 124
        4008 => X"71",  -- 113
        4009 => X"6A",  -- 106
        4010 => X"65",  -- 101
        4011 => X"68",  -- 104
        4012 => X"6F",  -- 111
        4013 => X"72",  -- 114
        4014 => X"71",  -- 113
        4015 => X"6C",  -- 108
        4016 => X"68",  -- 104
        4017 => X"6E",  -- 110
        4018 => X"75",  -- 117
        4019 => X"7B",  -- 123
        4020 => X"7E",  -- 126
        4021 => X"7F",  -- 127
        4022 => X"7D",  -- 125
        4023 => X"7C",  -- 124
        4024 => X"83",  -- 131
        4025 => X"7B",  -- 123
        4026 => X"83",  -- 131
        4027 => X"89",  -- 137
        4028 => X"83",  -- 131
        4029 => X"89",  -- 137
        4030 => X"8F",  -- 143
        4031 => X"86",  -- 134
        4032 => X"8C",  -- 140
        4033 => X"8D",  -- 141
        4034 => X"90",  -- 144
        4035 => X"91",  -- 145
        4036 => X"92",  -- 146
        4037 => X"93",  -- 147
        4038 => X"95",  -- 149
        4039 => X"95",  -- 149
        4040 => X"96",  -- 150
        4041 => X"9A",  -- 154
        4042 => X"9F",  -- 159
        4043 => X"A1",  -- 161
        4044 => X"A1",  -- 161
        4045 => X"A2",  -- 162
        4046 => X"A5",  -- 165
        4047 => X"A9",  -- 169
        4048 => X"A8",  -- 168
        4049 => X"AD",  -- 173
        4050 => X"B1",  -- 177
        4051 => X"B2",  -- 178
        4052 => X"B1",  -- 177
        4053 => X"B3",  -- 179
        4054 => X"B6",  -- 182
        4055 => X"BA",  -- 186
        4056 => X"BA",  -- 186
        4057 => X"B9",  -- 185
        4058 => X"B6",  -- 182
        4059 => X"B1",  -- 177
        4060 => X"B0",  -- 176
        4061 => X"AE",  -- 174
        4062 => X"A6",  -- 166
        4063 => X"9C",  -- 156
        4064 => X"99",  -- 153
        4065 => X"95",  -- 149
        4066 => X"94",  -- 148
        4067 => X"93",  -- 147
        4068 => X"90",  -- 144
        4069 => X"8D",  -- 141
        4070 => X"8F",  -- 143
        4071 => X"93",  -- 147
        4072 => X"9A",  -- 154
        4073 => X"9E",  -- 158
        4074 => X"A1",  -- 161
        4075 => X"A1",  -- 161
        4076 => X"9F",  -- 159
        4077 => X"9E",  -- 158
        4078 => X"A0",  -- 160
        4079 => X"A3",  -- 163
        4080 => X"9E",  -- 158
        4081 => X"9F",  -- 159
        4082 => X"A2",  -- 162
        4083 => X"A5",  -- 165
        4084 => X"A8",  -- 168
        4085 => X"A9",  -- 169
        4086 => X"A9",  -- 169
        4087 => X"A8",  -- 168
        4088 => X"AB",  -- 171
        4089 => X"A7",  -- 167
        4090 => X"AB",  -- 171
        4091 => X"B3",  -- 179
        4092 => X"B6",  -- 182
        4093 => X"B3",  -- 179
        4094 => X"B4",  -- 180
        4095 => X"BA",  -- 186
        4096 => X"B9",  -- 185
        4097 => X"B6",  -- 182
        4098 => X"B0",  -- 176
        4099 => X"AB",  -- 171
        4100 => X"A6",  -- 166
        4101 => X"A3",  -- 163
        4102 => X"9F",  -- 159
        4103 => X"9D",  -- 157
        4104 => X"9C",  -- 156
        4105 => X"9D",  -- 157
        4106 => X"9B",  -- 155
        4107 => X"97",  -- 151
        4108 => X"96",  -- 150
        4109 => X"93",  -- 147
        4110 => X"8B",  -- 139
        4111 => X"83",  -- 131
        4112 => X"8B",  -- 139
        4113 => X"85",  -- 133
        4114 => X"7D",  -- 125
        4115 => X"6E",  -- 110
        4116 => X"65",  -- 101
        4117 => X"6B",  -- 107
        4118 => X"65",  -- 101
        4119 => X"51",  -- 81
        4120 => X"44",  -- 68
        4121 => X"55",  -- 85
        4122 => X"68",  -- 104
        4123 => X"6E",  -- 110
        4124 => X"63",  -- 99
        4125 => X"57",  -- 87
        4126 => X"54",  -- 84
        4127 => X"56",  -- 86
        4128 => X"6F",  -- 111
        4129 => X"81",  -- 129
        4130 => X"93",  -- 147
        4131 => X"9D",  -- 157
        4132 => X"A6",  -- 166
        4133 => X"AF",  -- 175
        4134 => X"B5",  -- 181
        4135 => X"B2",  -- 178
        4136 => X"B6",  -- 182
        4137 => X"BA",  -- 186
        4138 => X"BE",  -- 190
        4139 => X"C2",  -- 194
        4140 => X"C2",  -- 194
        4141 => X"C2",  -- 194
        4142 => X"BF",  -- 191
        4143 => X"BF",  -- 191
        4144 => X"BF",  -- 191
        4145 => X"BC",  -- 188
        4146 => X"B8",  -- 184
        4147 => X"B5",  -- 181
        4148 => X"B4",  -- 180
        4149 => X"B3",  -- 179
        4150 => X"B4",  -- 180
        4151 => X"B6",  -- 182
        4152 => X"B8",  -- 184
        4153 => X"B7",  -- 183
        4154 => X"B6",  -- 182
        4155 => X"B6",  -- 182
        4156 => X"B3",  -- 179
        4157 => X"B0",  -- 176
        4158 => X"B1",  -- 177
        4159 => X"B7",  -- 183
        4160 => X"43",  -- 67
        4161 => X"41",  -- 65
        4162 => X"3F",  -- 63
        4163 => X"3D",  -- 61
        4164 => X"3B",  -- 59
        4165 => X"3A",  -- 58
        4166 => X"3A",  -- 58
        4167 => X"3B",  -- 59
        4168 => X"3B",  -- 59
        4169 => X"3A",  -- 58
        4170 => X"3A",  -- 58
        4171 => X"3A",  -- 58
        4172 => X"3B",  -- 59
        4173 => X"3C",  -- 60
        4174 => X"3E",  -- 62
        4175 => X"3E",  -- 62
        4176 => X"3E",  -- 62
        4177 => X"3E",  -- 62
        4178 => X"3E",  -- 62
        4179 => X"3E",  -- 62
        4180 => X"3E",  -- 62
        4181 => X"3E",  -- 62
        4182 => X"3E",  -- 62
        4183 => X"3E",  -- 62
        4184 => X"3E",  -- 62
        4185 => X"3E",  -- 62
        4186 => X"3F",  -- 63
        4187 => X"40",  -- 64
        4188 => X"40",  -- 64
        4189 => X"40",  -- 64
        4190 => X"3F",  -- 63
        4191 => X"3F",  -- 63
        4192 => X"3E",  -- 62
        4193 => X"3D",  -- 61
        4194 => X"3C",  -- 60
        4195 => X"3B",  -- 59
        4196 => X"3B",  -- 59
        4197 => X"3A",  -- 58
        4198 => X"39",  -- 57
        4199 => X"38",  -- 56
        4200 => X"38",  -- 56
        4201 => X"37",  -- 55
        4202 => X"35",  -- 53
        4203 => X"34",  -- 52
        4204 => X"33",  -- 51
        4205 => X"32",  -- 50
        4206 => X"31",  -- 49
        4207 => X"31",  -- 49
        4208 => X"30",  -- 48
        4209 => X"30",  -- 48
        4210 => X"30",  -- 48
        4211 => X"2F",  -- 47
        4212 => X"2E",  -- 46
        4213 => X"2C",  -- 44
        4214 => X"2B",  -- 43
        4215 => X"2A",  -- 42
        4216 => X"2A",  -- 42
        4217 => X"29",  -- 41
        4218 => X"28",  -- 40
        4219 => X"27",  -- 39
        4220 => X"27",  -- 39
        4221 => X"27",  -- 39
        4222 => X"28",  -- 40
        4223 => X"29",  -- 41
        4224 => X"2A",  -- 42
        4225 => X"2D",  -- 45
        4226 => X"30",  -- 48
        4227 => X"32",  -- 50
        4228 => X"35",  -- 53
        4229 => X"37",  -- 55
        4230 => X"3B",  -- 59
        4231 => X"3E",  -- 62
        4232 => X"3F",  -- 63
        4233 => X"40",  -- 64
        4234 => X"42",  -- 66
        4235 => X"45",  -- 69
        4236 => X"47",  -- 71
        4237 => X"49",  -- 73
        4238 => X"4A",  -- 74
        4239 => X"4A",  -- 74
        4240 => X"4E",  -- 78
        4241 => X"4D",  -- 77
        4242 => X"4B",  -- 75
        4243 => X"4A",  -- 74
        4244 => X"57",  -- 87
        4245 => X"73",  -- 115
        4246 => X"8F",  -- 143
        4247 => X"A2",  -- 162
        4248 => X"AA",  -- 170
        4249 => X"A1",  -- 161
        4250 => X"9C",  -- 156
        4251 => X"9D",  -- 157
        4252 => X"A2",  -- 162
        4253 => X"A4",  -- 164
        4254 => X"A1",  -- 161
        4255 => X"9C",  -- 156
        4256 => X"95",  -- 149
        4257 => X"98",  -- 152
        4258 => X"99",  -- 153
        4259 => X"99",  -- 153
        4260 => X"9C",  -- 156
        4261 => X"9C",  -- 156
        4262 => X"95",  -- 149
        4263 => X"8D",  -- 141
        4264 => X"8B",  -- 139
        4265 => X"82",  -- 130
        4266 => X"82",  -- 130
        4267 => X"75",  -- 117
        4268 => X"6E",  -- 110
        4269 => X"5C",  -- 92
        4270 => X"4E",  -- 78
        4271 => X"37",  -- 55
        4272 => X"36",  -- 54
        4273 => X"46",  -- 70
        4274 => X"71",  -- 113
        4275 => X"7A",  -- 122
        4276 => X"73",  -- 115
        4277 => X"74",  -- 116
        4278 => X"6F",  -- 111
        4279 => X"87",  -- 135
        4280 => X"86",  -- 134
        4281 => X"91",  -- 145
        4282 => X"89",  -- 137
        4283 => X"94",  -- 148
        4284 => X"99",  -- 153
        4285 => X"8C",  -- 140
        4286 => X"9C",  -- 156
        4287 => X"90",  -- 144
        4288 => X"95",  -- 149
        4289 => X"90",  -- 144
        4290 => X"8B",  -- 139
        4291 => X"89",  -- 137
        4292 => X"85",  -- 133
        4293 => X"7F",  -- 127
        4294 => X"7D",  -- 125
        4295 => X"7E",  -- 126
        4296 => X"72",  -- 114
        4297 => X"64",  -- 100
        4298 => X"61",  -- 97
        4299 => X"66",  -- 102
        4300 => X"64",  -- 100
        4301 => X"5C",  -- 92
        4302 => X"55",  -- 85
        4303 => X"4B",  -- 75
        4304 => X"4E",  -- 78
        4305 => X"45",  -- 69
        4306 => X"45",  -- 69
        4307 => X"51",  -- 81
        4308 => X"56",  -- 86
        4309 => X"50",  -- 80
        4310 => X"4F",  -- 79
        4311 => X"53",  -- 83
        4312 => X"56",  -- 86
        4313 => X"61",  -- 97
        4314 => X"6C",  -- 108
        4315 => X"72",  -- 114
        4316 => X"7D",  -- 125
        4317 => X"8A",  -- 138
        4318 => X"93",  -- 147
        4319 => X"94",  -- 148
        4320 => X"9D",  -- 157
        4321 => X"A3",  -- 163
        4322 => X"A8",  -- 168
        4323 => X"A9",  -- 169
        4324 => X"A1",  -- 161
        4325 => X"8D",  -- 141
        4326 => X"77",  -- 119
        4327 => X"68",  -- 104
        4328 => X"6D",  -- 109
        4329 => X"63",  -- 99
        4330 => X"5F",  -- 95
        4331 => X"63",  -- 99
        4332 => X"6D",  -- 109
        4333 => X"70",  -- 112
        4334 => X"6F",  -- 111
        4335 => X"6F",  -- 111
        4336 => X"72",  -- 114
        4337 => X"77",  -- 119
        4338 => X"78",  -- 120
        4339 => X"75",  -- 117
        4340 => X"74",  -- 116
        4341 => X"77",  -- 119
        4342 => X"7A",  -- 122
        4343 => X"7C",  -- 124
        4344 => X"82",  -- 130
        4345 => X"7F",  -- 127
        4346 => X"84",  -- 132
        4347 => X"89",  -- 137
        4348 => X"87",  -- 135
        4349 => X"89",  -- 137
        4350 => X"89",  -- 137
        4351 => X"83",  -- 131
        4352 => X"88",  -- 136
        4353 => X"8A",  -- 138
        4354 => X"8E",  -- 142
        4355 => X"90",  -- 144
        4356 => X"91",  -- 145
        4357 => X"92",  -- 146
        4358 => X"94",  -- 148
        4359 => X"95",  -- 149
        4360 => X"91",  -- 145
        4361 => X"95",  -- 149
        4362 => X"9A",  -- 154
        4363 => X"9C",  -- 156
        4364 => X"9C",  -- 156
        4365 => X"9D",  -- 157
        4366 => X"A2",  -- 162
        4367 => X"A7",  -- 167
        4368 => X"A8",  -- 168
        4369 => X"AE",  -- 174
        4370 => X"B4",  -- 180
        4371 => X"B4",  -- 180
        4372 => X"B1",  -- 177
        4373 => X"B2",  -- 178
        4374 => X"B5",  -- 181
        4375 => X"B9",  -- 185
        4376 => X"B8",  -- 184
        4377 => X"BA",  -- 186
        4378 => X"BA",  -- 186
        4379 => X"B4",  -- 180
        4380 => X"B1",  -- 177
        4381 => X"AD",  -- 173
        4382 => X"A5",  -- 165
        4383 => X"9C",  -- 156
        4384 => X"92",  -- 146
        4385 => X"8F",  -- 143
        4386 => X"8F",  -- 143
        4387 => X"90",  -- 144
        4388 => X"8F",  -- 143
        4389 => X"8D",  -- 141
        4390 => X"90",  -- 144
        4391 => X"95",  -- 149
        4392 => X"9E",  -- 158
        4393 => X"A2",  -- 162
        4394 => X"A4",  -- 164
        4395 => X"A2",  -- 162
        4396 => X"9E",  -- 158
        4397 => X"9C",  -- 156
        4398 => X"9F",  -- 159
        4399 => X"A3",  -- 163
        4400 => X"A1",  -- 161
        4401 => X"A1",  -- 161
        4402 => X"A3",  -- 163
        4403 => X"A6",  -- 166
        4404 => X"A9",  -- 169
        4405 => X"AA",  -- 170
        4406 => X"A7",  -- 167
        4407 => X"A4",  -- 164
        4408 => X"AC",  -- 172
        4409 => X"AC",  -- 172
        4410 => X"B1",  -- 177
        4411 => X"B7",  -- 183
        4412 => X"B9",  -- 185
        4413 => X"B7",  -- 183
        4414 => X"B5",  -- 181
        4415 => X"B8",  -- 184
        4416 => X"B6",  -- 182
        4417 => X"B6",  -- 182
        4418 => X"B4",  -- 180
        4419 => X"B1",  -- 177
        4420 => X"AD",  -- 173
        4421 => X"A7",  -- 167
        4422 => X"A1",  -- 161
        4423 => X"9F",  -- 159
        4424 => X"A1",  -- 161
        4425 => X"A3",  -- 163
        4426 => X"A2",  -- 162
        4427 => X"9D",  -- 157
        4428 => X"98",  -- 152
        4429 => X"97",  -- 151
        4430 => X"93",  -- 147
        4431 => X"90",  -- 144
        4432 => X"88",  -- 136
        4433 => X"85",  -- 133
        4434 => X"85",  -- 133
        4435 => X"82",  -- 130
        4436 => X"7F",  -- 127
        4437 => X"82",  -- 130
        4438 => X"75",  -- 117
        4439 => X"5D",  -- 93
        4440 => X"4B",  -- 75
        4441 => X"57",  -- 87
        4442 => X"60",  -- 96
        4443 => X"5F",  -- 95
        4444 => X"59",  -- 89
        4445 => X"56",  -- 86
        4446 => X"58",  -- 88
        4447 => X"59",  -- 89
        4448 => X"63",  -- 99
        4449 => X"6F",  -- 111
        4450 => X"7F",  -- 127
        4451 => X"8A",  -- 138
        4452 => X"95",  -- 149
        4453 => X"A2",  -- 162
        4454 => X"B0",  -- 176
        4455 => X"B6",  -- 182
        4456 => X"BE",  -- 190
        4457 => X"BE",  -- 190
        4458 => X"BD",  -- 189
        4459 => X"BE",  -- 190
        4460 => X"BD",  -- 189
        4461 => X"BD",  -- 189
        4462 => X"BF",  -- 191
        4463 => X"C1",  -- 193
        4464 => X"C5",  -- 197
        4465 => X"C1",  -- 193
        4466 => X"BF",  -- 191
        4467 => X"BF",  -- 191
        4468 => X"BD",  -- 189
        4469 => X"B9",  -- 185
        4470 => X"B7",  -- 183
        4471 => X"B8",  -- 184
        4472 => X"B6",  -- 182
        4473 => X"B3",  -- 179
        4474 => X"B1",  -- 177
        4475 => X"B2",  -- 178
        4476 => X"B2",  -- 178
        4477 => X"B2",  -- 178
        4478 => X"B5",  -- 181
        4479 => X"BB",  -- 187
        4480 => X"43",  -- 67
        4481 => X"41",  -- 65
        4482 => X"3F",  -- 63
        4483 => X"3D",  -- 61
        4484 => X"3A",  -- 58
        4485 => X"3A",  -- 58
        4486 => X"3A",  -- 58
        4487 => X"3A",  -- 58
        4488 => X"3B",  -- 59
        4489 => X"3B",  -- 59
        4490 => X"3A",  -- 58
        4491 => X"3B",  -- 59
        4492 => X"3B",  -- 59
        4493 => X"3C",  -- 60
        4494 => X"3E",  -- 62
        4495 => X"3F",  -- 63
        4496 => X"3F",  -- 63
        4497 => X"3F",  -- 63
        4498 => X"3F",  -- 63
        4499 => X"3F",  -- 63
        4500 => X"3F",  -- 63
        4501 => X"3F",  -- 63
        4502 => X"3F",  -- 63
        4503 => X"3F",  -- 63
        4504 => X"3E",  -- 62
        4505 => X"3E",  -- 62
        4506 => X"3F",  -- 63
        4507 => X"40",  -- 64
        4508 => X"40",  -- 64
        4509 => X"40",  -- 64
        4510 => X"40",  -- 64
        4511 => X"3F",  -- 63
        4512 => X"3E",  -- 62
        4513 => X"3E",  -- 62
        4514 => X"3D",  -- 61
        4515 => X"3B",  -- 59
        4516 => X"3B",  -- 59
        4517 => X"3A",  -- 58
        4518 => X"39",  -- 57
        4519 => X"38",  -- 56
        4520 => X"38",  -- 56
        4521 => X"37",  -- 55
        4522 => X"36",  -- 54
        4523 => X"35",  -- 53
        4524 => X"33",  -- 51
        4525 => X"32",  -- 50
        4526 => X"32",  -- 50
        4527 => X"31",  -- 49
        4528 => X"30",  -- 48
        4529 => X"30",  -- 48
        4530 => X"30",  -- 48
        4531 => X"2F",  -- 47
        4532 => X"2E",  -- 46
        4533 => X"2D",  -- 45
        4534 => X"2B",  -- 43
        4535 => X"2B",  -- 43
        4536 => X"2B",  -- 43
        4537 => X"2A",  -- 42
        4538 => X"29",  -- 41
        4539 => X"28",  -- 40
        4540 => X"27",  -- 39
        4541 => X"28",  -- 40
        4542 => X"29",  -- 41
        4543 => X"29",  -- 41
        4544 => X"2A",  -- 42
        4545 => X"2D",  -- 45
        4546 => X"30",  -- 48
        4547 => X"33",  -- 51
        4548 => X"35",  -- 53
        4549 => X"38",  -- 56
        4550 => X"3C",  -- 60
        4551 => X"3F",  -- 63
        4552 => X"40",  -- 64
        4553 => X"41",  -- 65
        4554 => X"43",  -- 67
        4555 => X"46",  -- 70
        4556 => X"48",  -- 72
        4557 => X"49",  -- 73
        4558 => X"4A",  -- 74
        4559 => X"4B",  -- 75
        4560 => X"4D",  -- 77
        4561 => X"50",  -- 80
        4562 => X"52",  -- 82
        4563 => X"58",  -- 88
        4564 => X"69",  -- 105
        4565 => X"85",  -- 133
        4566 => X"9E",  -- 158
        4567 => X"AB",  -- 171
        4568 => X"A6",  -- 166
        4569 => X"A0",  -- 160
        4570 => X"9B",  -- 155
        4571 => X"99",  -- 153
        4572 => X"9F",  -- 159
        4573 => X"A4",  -- 164
        4574 => X"A2",  -- 162
        4575 => X"9E",  -- 158
        4576 => X"95",  -- 149
        4577 => X"9A",  -- 154
        4578 => X"99",  -- 153
        4579 => X"97",  -- 151
        4580 => X"9C",  -- 156
        4581 => X"9A",  -- 154
        4582 => X"90",  -- 144
        4583 => X"8B",  -- 139
        4584 => X"89",  -- 137
        4585 => X"7C",  -- 124
        4586 => X"7D",  -- 125
        4587 => X"6D",  -- 109
        4588 => X"63",  -- 99
        4589 => X"4B",  -- 75
        4590 => X"47",  -- 71
        4591 => X"39",  -- 57
        4592 => X"46",  -- 70
        4593 => X"59",  -- 89
        4594 => X"74",  -- 116
        4595 => X"82",  -- 130
        4596 => X"83",  -- 131
        4597 => X"7E",  -- 126
        4598 => X"7F",  -- 127
        4599 => X"87",  -- 135
        4600 => X"8E",  -- 142
        4601 => X"8F",  -- 143
        4602 => X"8B",  -- 139
        4603 => X"96",  -- 150
        4604 => X"93",  -- 147
        4605 => X"91",  -- 145
        4606 => X"90",  -- 144
        4607 => X"93",  -- 147
        4608 => X"90",  -- 144
        4609 => X"8E",  -- 142
        4610 => X"8A",  -- 138
        4611 => X"82",  -- 130
        4612 => X"7D",  -- 125
        4613 => X"77",  -- 119
        4614 => X"72",  -- 114
        4615 => X"6C",  -- 108
        4616 => X"62",  -- 98
        4617 => X"58",  -- 88
        4618 => X"52",  -- 82
        4619 => X"5A",  -- 90
        4620 => X"5E",  -- 94
        4621 => X"4E",  -- 78
        4622 => X"3F",  -- 63
        4623 => X"41",  -- 65
        4624 => X"42",  -- 66
        4625 => X"3F",  -- 63
        4626 => X"41",  -- 65
        4627 => X"45",  -- 69
        4628 => X"42",  -- 66
        4629 => X"3C",  -- 60
        4630 => X"40",  -- 64
        4631 => X"4B",  -- 75
        4632 => X"52",  -- 82
        4633 => X"55",  -- 85
        4634 => X"5A",  -- 90
        4635 => X"5D",  -- 93
        4636 => X"62",  -- 98
        4637 => X"72",  -- 114
        4638 => X"84",  -- 132
        4639 => X"93",  -- 147
        4640 => X"AE",  -- 174
        4641 => X"AA",  -- 170
        4642 => X"A2",  -- 162
        4643 => X"9B",  -- 155
        4644 => X"94",  -- 148
        4645 => X"86",  -- 134
        4646 => X"78",  -- 120
        4647 => X"6E",  -- 110
        4648 => X"62",  -- 98
        4649 => X"5E",  -- 94
        4650 => X"5D",  -- 93
        4651 => X"61",  -- 97
        4652 => X"67",  -- 103
        4653 => X"6B",  -- 107
        4654 => X"6E",  -- 110
        4655 => X"72",  -- 114
        4656 => X"77",  -- 119
        4657 => X"79",  -- 121
        4658 => X"78",  -- 120
        4659 => X"71",  -- 113
        4660 => X"6D",  -- 109
        4661 => X"73",  -- 115
        4662 => X"7B",  -- 123
        4663 => X"7F",  -- 127
        4664 => X"80",  -- 128
        4665 => X"84",  -- 132
        4666 => X"83",  -- 131
        4667 => X"83",  -- 131
        4668 => X"88",  -- 136
        4669 => X"85",  -- 133
        4670 => X"7E",  -- 126
        4671 => X"7F",  -- 127
        4672 => X"7E",  -- 126
        4673 => X"83",  -- 131
        4674 => X"88",  -- 136
        4675 => X"8D",  -- 141
        4676 => X"90",  -- 144
        4677 => X"92",  -- 146
        4678 => X"95",  -- 149
        4679 => X"97",  -- 151
        4680 => X"91",  -- 145
        4681 => X"95",  -- 149
        4682 => X"99",  -- 153
        4683 => X"99",  -- 153
        4684 => X"98",  -- 152
        4685 => X"99",  -- 153
        4686 => X"A0",  -- 160
        4687 => X"A5",  -- 165
        4688 => X"AA",  -- 170
        4689 => X"AE",  -- 174
        4690 => X"B2",  -- 178
        4691 => X"B4",  -- 180
        4692 => X"B2",  -- 178
        4693 => X"B3",  -- 179
        4694 => X"B3",  -- 179
        4695 => X"B4",  -- 180
        4696 => X"B5",  -- 181
        4697 => X"BA",  -- 186
        4698 => X"BE",  -- 190
        4699 => X"B8",  -- 184
        4700 => X"B2",  -- 178
        4701 => X"AB",  -- 171
        4702 => X"A4",  -- 164
        4703 => X"9C",  -- 156
        4704 => X"8E",  -- 142
        4705 => X"8B",  -- 139
        4706 => X"8A",  -- 138
        4707 => X"8D",  -- 141
        4708 => X"8F",  -- 143
        4709 => X"90",  -- 144
        4710 => X"97",  -- 151
        4711 => X"9E",  -- 158
        4712 => X"9F",  -- 159
        4713 => X"A0",  -- 160
        4714 => X"A0",  -- 160
        4715 => X"9F",  -- 159
        4716 => X"9D",  -- 157
        4717 => X"9D",  -- 157
        4718 => X"A0",  -- 160
        4719 => X"A3",  -- 163
        4720 => X"A3",  -- 163
        4721 => X"A4",  -- 164
        4722 => X"A5",  -- 165
        4723 => X"A6",  -- 166
        4724 => X"A6",  -- 166
        4725 => X"A6",  -- 166
        4726 => X"A7",  -- 167
        4727 => X"A7",  -- 167
        4728 => X"AD",  -- 173
        4729 => X"B2",  -- 178
        4730 => X"B6",  -- 182
        4731 => X"B6",  -- 182
        4732 => X"B7",  -- 183
        4733 => X"B9",  -- 185
        4734 => X"B6",  -- 182
        4735 => X"B4",  -- 180
        4736 => X"B5",  -- 181
        4737 => X"B6",  -- 182
        4738 => X"B7",  -- 183
        4739 => X"B5",  -- 181
        4740 => X"AF",  -- 175
        4741 => X"AA",  -- 170
        4742 => X"A4",  -- 164
        4743 => X"A1",  -- 161
        4744 => X"A1",  -- 161
        4745 => X"A4",  -- 164
        4746 => X"A2",  -- 162
        4747 => X"9C",  -- 156
        4748 => X"98",  -- 152
        4749 => X"98",  -- 152
        4750 => X"99",  -- 153
        4751 => X"96",  -- 150
        4752 => X"8D",  -- 141
        4753 => X"8B",  -- 139
        4754 => X"92",  -- 146
        4755 => X"96",  -- 150
        4756 => X"94",  -- 148
        4757 => X"92",  -- 146
        4758 => X"84",  -- 132
        4759 => X"6E",  -- 110
        4760 => X"60",  -- 96
        4761 => X"62",  -- 98
        4762 => X"60",  -- 96
        4763 => X"5F",  -- 95
        4764 => X"60",  -- 96
        4765 => X"63",  -- 99
        4766 => X"5E",  -- 94
        4767 => X"55",  -- 85
        4768 => X"53",  -- 83
        4769 => X"5E",  -- 94
        4770 => X"6C",  -- 108
        4771 => X"76",  -- 118
        4772 => X"7C",  -- 124
        4773 => X"88",  -- 136
        4774 => X"A1",  -- 161
        4775 => X"B8",  -- 184
        4776 => X"BB",  -- 187
        4777 => X"BB",  -- 187
        4778 => X"BA",  -- 186
        4779 => X"BB",  -- 187
        4780 => X"BB",  -- 187
        4781 => X"BC",  -- 188
        4782 => X"C0",  -- 192
        4783 => X"C2",  -- 194
        4784 => X"C5",  -- 197
        4785 => X"C2",  -- 194
        4786 => X"C2",  -- 194
        4787 => X"C5",  -- 197
        4788 => X"C3",  -- 195
        4789 => X"BC",  -- 188
        4790 => X"B7",  -- 183
        4791 => X"B7",  -- 183
        4792 => X"B6",  -- 182
        4793 => X"B1",  -- 177
        4794 => X"AF",  -- 175
        4795 => X"B2",  -- 178
        4796 => X"B4",  -- 180
        4797 => X"B5",  -- 181
        4798 => X"B7",  -- 183
        4799 => X"BB",  -- 187
        4800 => X"43",  -- 67
        4801 => X"41",  -- 65
        4802 => X"3F",  -- 63
        4803 => X"3D",  -- 61
        4804 => X"3A",  -- 58
        4805 => X"39",  -- 57
        4806 => X"39",  -- 57
        4807 => X"3A",  -- 58
        4808 => X"3B",  -- 59
        4809 => X"3B",  -- 59
        4810 => X"3B",  -- 59
        4811 => X"3B",  -- 59
        4812 => X"3B",  -- 59
        4813 => X"3C",  -- 60
        4814 => X"3D",  -- 61
        4815 => X"3E",  -- 62
        4816 => X"3F",  -- 63
        4817 => X"3F",  -- 63
        4818 => X"3F",  -- 63
        4819 => X"3F",  -- 63
        4820 => X"3F",  -- 63
        4821 => X"3F",  -- 63
        4822 => X"3F",  -- 63
        4823 => X"3F",  -- 63
        4824 => X"3E",  -- 62
        4825 => X"3F",  -- 63
        4826 => X"3F",  -- 63
        4827 => X"40",  -- 64
        4828 => X"40",  -- 64
        4829 => X"40",  -- 64
        4830 => X"40",  -- 64
        4831 => X"3F",  -- 63
        4832 => X"3E",  -- 62
        4833 => X"3E",  -- 62
        4834 => X"3D",  -- 61
        4835 => X"3C",  -- 60
        4836 => X"3B",  -- 59
        4837 => X"3A",  -- 58
        4838 => X"39",  -- 57
        4839 => X"38",  -- 56
        4840 => X"38",  -- 56
        4841 => X"36",  -- 54
        4842 => X"36",  -- 54
        4843 => X"35",  -- 53
        4844 => X"34",  -- 52
        4845 => X"33",  -- 51
        4846 => X"32",  -- 50
        4847 => X"31",  -- 49
        4848 => X"31",  -- 49
        4849 => X"31",  -- 49
        4850 => X"31",  -- 49
        4851 => X"30",  -- 48
        4852 => X"2F",  -- 47
        4853 => X"2D",  -- 45
        4854 => X"2C",  -- 44
        4855 => X"2B",  -- 43
        4856 => X"2B",  -- 43
        4857 => X"2A",  -- 42
        4858 => X"29",  -- 41
        4859 => X"28",  -- 40
        4860 => X"28",  -- 40
        4861 => X"28",  -- 40
        4862 => X"29",  -- 41
        4863 => X"2A",  -- 42
        4864 => X"2B",  -- 43
        4865 => X"2E",  -- 46
        4866 => X"31",  -- 49
        4867 => X"33",  -- 51
        4868 => X"35",  -- 53
        4869 => X"39",  -- 57
        4870 => X"3C",  -- 60
        4871 => X"3E",  -- 62
        4872 => X"40",  -- 64
        4873 => X"41",  -- 65
        4874 => X"43",  -- 67
        4875 => X"46",  -- 70
        4876 => X"48",  -- 72
        4877 => X"4B",  -- 75
        4878 => X"4B",  -- 75
        4879 => X"4C",  -- 76
        4880 => X"48",  -- 72
        4881 => X"52",  -- 82
        4882 => X"5D",  -- 93
        4883 => X"6A",  -- 106
        4884 => X"7E",  -- 126
        4885 => X"94",  -- 148
        4886 => X"A4",  -- 164
        4887 => X"A8",  -- 168
        4888 => X"A5",  -- 165
        4889 => X"A3",  -- 163
        4890 => X"9E",  -- 158
        4891 => X"9B",  -- 155
        4892 => X"A0",  -- 160
        4893 => X"A5",  -- 165
        4894 => X"A7",  -- 167
        4895 => X"A2",  -- 162
        4896 => X"90",  -- 144
        4897 => X"9A",  -- 154
        4898 => X"9C",  -- 156
        4899 => X"9B",  -- 155
        4900 => X"9E",  -- 158
        4901 => X"97",  -- 151
        4902 => X"8B",  -- 139
        4903 => X"85",  -- 133
        4904 => X"88",  -- 136
        4905 => X"76",  -- 118
        4906 => X"78",  -- 120
        4907 => X"66",  -- 102
        4908 => X"5B",  -- 91
        4909 => X"3F",  -- 63
        4910 => X"41",  -- 65
        4911 => X"3B",  -- 59
        4912 => X"58",  -- 88
        4913 => X"68",  -- 104
        4914 => X"71",  -- 113
        4915 => X"81",  -- 129
        4916 => X"84",  -- 132
        4917 => X"84",  -- 132
        4918 => X"8C",  -- 140
        4919 => X"8E",  -- 142
        4920 => X"95",  -- 149
        4921 => X"89",  -- 137
        4922 => X"8F",  -- 143
        4923 => X"98",  -- 152
        4924 => X"8C",  -- 140
        4925 => X"96",  -- 150
        4926 => X"83",  -- 131
        4927 => X"97",  -- 151
        4928 => X"8E",  -- 142
        4929 => X"90",  -- 144
        4930 => X"8D",  -- 141
        4931 => X"80",  -- 128
        4932 => X"78",  -- 120
        4933 => X"71",  -- 113
        4934 => X"67",  -- 103
        4935 => X"5D",  -- 93
        4936 => X"5B",  -- 91
        4937 => X"5A",  -- 90
        4938 => X"49",  -- 73
        4939 => X"44",  -- 68
        4940 => X"55",  -- 85
        4941 => X"53",  -- 83
        4942 => X"40",  -- 64
        4943 => X"39",  -- 57
        4944 => X"35",  -- 53
        4945 => X"34",  -- 52
        4946 => X"35",  -- 53
        4947 => X"38",  -- 56
        4948 => X"3B",  -- 59
        4949 => X"42",  -- 66
        4950 => X"4E",  -- 78
        4951 => X"58",  -- 88
        4952 => X"48",  -- 72
        4953 => X"49",  -- 73
        4954 => X"4B",  -- 75
        4955 => X"4C",  -- 76
        4956 => X"52",  -- 82
        4957 => X"64",  -- 100
        4958 => X"83",  -- 131
        4959 => X"9D",  -- 157
        4960 => X"A1",  -- 161
        4961 => X"9F",  -- 159
        4962 => X"9D",  -- 157
        4963 => X"9A",  -- 154
        4964 => X"96",  -- 150
        4965 => X"8B",  -- 139
        4966 => X"78",  -- 120
        4967 => X"6B",  -- 107
        4968 => X"5D",  -- 93
        4969 => X"5B",  -- 91
        4970 => X"5C",  -- 92
        4971 => X"60",  -- 96
        4972 => X"62",  -- 98
        4973 => X"63",  -- 99
        4974 => X"6A",  -- 106
        4975 => X"72",  -- 114
        4976 => X"72",  -- 114
        4977 => X"77",  -- 119
        4978 => X"76",  -- 118
        4979 => X"70",  -- 112
        4980 => X"6C",  -- 108
        4981 => X"74",  -- 116
        4982 => X"7B",  -- 123
        4983 => X"80",  -- 128
        4984 => X"7D",  -- 125
        4985 => X"85",  -- 133
        4986 => X"7E",  -- 126
        4987 => X"7C",  -- 124
        4988 => X"85",  -- 133
        4989 => X"80",  -- 128
        4990 => X"77",  -- 119
        4991 => X"7D",  -- 125
        4992 => X"7F",  -- 127
        4993 => X"83",  -- 131
        4994 => X"89",  -- 137
        4995 => X"8C",  -- 140
        4996 => X"8E",  -- 142
        4997 => X"8E",  -- 142
        4998 => X"90",  -- 144
        4999 => X"91",  -- 145
        5000 => X"93",  -- 147
        5001 => X"97",  -- 151
        5002 => X"9A",  -- 154
        5003 => X"99",  -- 153
        5004 => X"97",  -- 151
        5005 => X"99",  -- 153
        5006 => X"9F",  -- 159
        5007 => X"A4",  -- 164
        5008 => X"AC",  -- 172
        5009 => X"AD",  -- 173
        5010 => X"AF",  -- 175
        5011 => X"B2",  -- 178
        5012 => X"B4",  -- 180
        5013 => X"B5",  -- 181
        5014 => X"B2",  -- 178
        5015 => X"B0",  -- 176
        5016 => X"B3",  -- 179
        5017 => X"BB",  -- 187
        5018 => X"C0",  -- 192
        5019 => X"BC",  -- 188
        5020 => X"B1",  -- 177
        5021 => X"A9",  -- 169
        5022 => X"A3",  -- 163
        5023 => X"9C",  -- 156
        5024 => X"92",  -- 146
        5025 => X"8C",  -- 140
        5026 => X"89",  -- 137
        5027 => X"89",  -- 137
        5028 => X"8A",  -- 138
        5029 => X"8B",  -- 139
        5030 => X"92",  -- 146
        5031 => X"99",  -- 153
        5032 => X"9C",  -- 156
        5033 => X"9A",  -- 154
        5034 => X"99",  -- 153
        5035 => X"99",  -- 153
        5036 => X"9B",  -- 155
        5037 => X"9F",  -- 159
        5038 => X"A1",  -- 161
        5039 => X"A2",  -- 162
        5040 => X"A3",  -- 163
        5041 => X"A5",  -- 165
        5042 => X"A7",  -- 167
        5043 => X"A5",  -- 165
        5044 => X"A2",  -- 162
        5045 => X"A3",  -- 163
        5046 => X"A9",  -- 169
        5047 => X"AE",  -- 174
        5048 => X"AE",  -- 174
        5049 => X"B4",  -- 180
        5050 => X"B7",  -- 183
        5051 => X"B3",  -- 179
        5052 => X"B3",  -- 179
        5053 => X"B8",  -- 184
        5054 => X"B6",  -- 182
        5055 => X"B1",  -- 177
        5056 => X"B5",  -- 181
        5057 => X"B6",  -- 182
        5058 => X"B6",  -- 182
        5059 => X"B4",  -- 180
        5060 => X"B0",  -- 176
        5061 => X"AB",  -- 171
        5062 => X"A7",  -- 167
        5063 => X"A3",  -- 163
        5064 => X"A0",  -- 160
        5065 => X"A0",  -- 160
        5066 => X"9D",  -- 157
        5067 => X"99",  -- 153
        5068 => X"96",  -- 150
        5069 => X"9A",  -- 154
        5070 => X"9A",  -- 154
        5071 => X"97",  -- 151
        5072 => X"99",  -- 153
        5073 => X"97",  -- 151
        5074 => X"9D",  -- 157
        5075 => X"A2",  -- 162
        5076 => X"9C",  -- 156
        5077 => X"95",  -- 149
        5078 => X"89",  -- 137
        5079 => X"78",  -- 120
        5080 => X"71",  -- 113
        5081 => X"6D",  -- 109
        5082 => X"66",  -- 102
        5083 => X"65",  -- 101
        5084 => X"6C",  -- 108
        5085 => X"6D",  -- 109
        5086 => X"5D",  -- 93
        5087 => X"48",  -- 72
        5088 => X"51",  -- 81
        5089 => X"59",  -- 89
        5090 => X"66",  -- 102
        5091 => X"69",  -- 105
        5092 => X"65",  -- 101
        5093 => X"6D",  -- 109
        5094 => X"8B",  -- 139
        5095 => X"AC",  -- 172
        5096 => X"B0",  -- 176
        5097 => X"B4",  -- 180
        5098 => X"B9",  -- 185
        5099 => X"BC",  -- 188
        5100 => X"BF",  -- 191
        5101 => X"C1",  -- 193
        5102 => X"C1",  -- 193
        5103 => X"C2",  -- 194
        5104 => X"BF",  -- 191
        5105 => X"BE",  -- 190
        5106 => X"C1",  -- 193
        5107 => X"C5",  -- 197
        5108 => X"C3",  -- 195
        5109 => X"BA",  -- 186
        5110 => X"B3",  -- 179
        5111 => X"B2",  -- 178
        5112 => X"BA",  -- 186
        5113 => X"B4",  -- 180
        5114 => X"B1",  -- 177
        5115 => X"B4",  -- 180
        5116 => X"B8",  -- 184
        5117 => X"B7",  -- 183
        5118 => X"B7",  -- 183
        5119 => X"B8",  -- 184
        5120 => X"3F",  -- 63
        5121 => X"3E",  -- 62
        5122 => X"3D",  -- 61
        5123 => X"3B",  -- 59
        5124 => X"3A",  -- 58
        5125 => X"3A",  -- 58
        5126 => X"3A",  -- 58
        5127 => X"3A",  -- 58
        5128 => X"3A",  -- 58
        5129 => X"3A",  -- 58
        5130 => X"3B",  -- 59
        5131 => X"3B",  -- 59
        5132 => X"3C",  -- 60
        5133 => X"3C",  -- 60
        5134 => X"3D",  -- 61
        5135 => X"3D",  -- 61
        5136 => X"3D",  -- 61
        5137 => X"3D",  -- 61
        5138 => X"3D",  -- 61
        5139 => X"3D",  -- 61
        5140 => X"3D",  -- 61
        5141 => X"3D",  -- 61
        5142 => X"3D",  -- 61
        5143 => X"3D",  -- 61
        5144 => X"3D",  -- 61
        5145 => X"3D",  -- 61
        5146 => X"3F",  -- 63
        5147 => X"40",  -- 64
        5148 => X"40",  -- 64
        5149 => X"41",  -- 65
        5150 => X"41",  -- 65
        5151 => X"41",  -- 65
        5152 => X"3E",  -- 62
        5153 => X"3E",  -- 62
        5154 => X"3D",  -- 61
        5155 => X"3C",  -- 60
        5156 => X"3A",  -- 58
        5157 => X"3A",  -- 58
        5158 => X"39",  -- 57
        5159 => X"38",  -- 56
        5160 => X"37",  -- 55
        5161 => X"35",  -- 53
        5162 => X"35",  -- 53
        5163 => X"34",  -- 52
        5164 => X"33",  -- 51
        5165 => X"33",  -- 51
        5166 => X"32",  -- 50
        5167 => X"32",  -- 50
        5168 => X"31",  -- 49
        5169 => X"30",  -- 48
        5170 => X"31",  -- 49
        5171 => X"30",  -- 48
        5172 => X"2F",  -- 47
        5173 => X"2D",  -- 45
        5174 => X"2D",  -- 45
        5175 => X"2D",  -- 45
        5176 => X"2B",  -- 43
        5177 => X"29",  -- 41
        5178 => X"27",  -- 39
        5179 => X"27",  -- 39
        5180 => X"28",  -- 40
        5181 => X"29",  -- 41
        5182 => X"2A",  -- 42
        5183 => X"28",  -- 40
        5184 => X"2D",  -- 45
        5185 => X"2F",  -- 47
        5186 => X"32",  -- 50
        5187 => X"34",  -- 52
        5188 => X"37",  -- 55
        5189 => X"39",  -- 57
        5190 => X"3E",  -- 62
        5191 => X"3F",  -- 63
        5192 => X"41",  -- 65
        5193 => X"44",  -- 68
        5194 => X"47",  -- 71
        5195 => X"47",  -- 71
        5196 => X"47",  -- 71
        5197 => X"49",  -- 73
        5198 => X"4E",  -- 78
        5199 => X"50",  -- 80
        5200 => X"4E",  -- 78
        5201 => X"5A",  -- 90
        5202 => X"69",  -- 105
        5203 => X"88",  -- 136
        5204 => X"94",  -- 148
        5205 => X"92",  -- 146
        5206 => X"A4",  -- 164
        5207 => X"B0",  -- 176
        5208 => X"A6",  -- 166
        5209 => X"A7",  -- 167
        5210 => X"A2",  -- 162
        5211 => X"9C",  -- 156
        5212 => X"9C",  -- 156
        5213 => X"A5",  -- 165
        5214 => X"A9",  -- 169
        5215 => X"A6",  -- 166
        5216 => X"96",  -- 150
        5217 => X"90",  -- 144
        5218 => X"9C",  -- 156
        5219 => X"A1",  -- 161
        5220 => X"9D",  -- 157
        5221 => X"95",  -- 149
        5222 => X"87",  -- 135
        5223 => X"8B",  -- 139
        5224 => X"81",  -- 129
        5225 => X"79",  -- 121
        5226 => X"74",  -- 116
        5227 => X"59",  -- 89
        5228 => X"4D",  -- 77
        5229 => X"3A",  -- 58
        5230 => X"43",  -- 67
        5231 => X"48",  -- 72
        5232 => X"5E",  -- 94
        5233 => X"66",  -- 102
        5234 => X"71",  -- 113
        5235 => X"87",  -- 135
        5236 => X"7A",  -- 122
        5237 => X"86",  -- 134
        5238 => X"8B",  -- 139
        5239 => X"94",  -- 148
        5240 => X"94",  -- 148
        5241 => X"8F",  -- 143
        5242 => X"8D",  -- 141
        5243 => X"90",  -- 144
        5244 => X"95",  -- 149
        5245 => X"98",  -- 152
        5246 => X"95",  -- 149
        5247 => X"93",  -- 147
        5248 => X"84",  -- 132
        5249 => X"8D",  -- 141
        5250 => X"95",  -- 149
        5251 => X"85",  -- 133
        5252 => X"6A",  -- 106
        5253 => X"67",  -- 103
        5254 => X"64",  -- 100
        5255 => X"4F",  -- 79
        5256 => X"52",  -- 82
        5257 => X"54",  -- 84
        5258 => X"4F",  -- 79
        5259 => X"50",  -- 80
        5260 => X"52",  -- 82
        5261 => X"3D",  -- 61
        5262 => X"31",  -- 49
        5263 => X"3E",  -- 62
        5264 => X"3C",  -- 60
        5265 => X"41",  -- 65
        5266 => X"40",  -- 64
        5267 => X"3F",  -- 63
        5268 => X"4D",  -- 77
        5269 => X"5E",  -- 94
        5270 => X"57",  -- 87
        5271 => X"43",  -- 67
        5272 => X"49",  -- 73
        5273 => X"46",  -- 70
        5274 => X"40",  -- 64
        5275 => X"41",  -- 65
        5276 => X"4E",  -- 78
        5277 => X"63",  -- 99
        5278 => X"73",  -- 115
        5279 => X"78",  -- 120
        5280 => X"86",  -- 134
        5281 => X"92",  -- 146
        5282 => X"99",  -- 153
        5283 => X"8F",  -- 143
        5284 => X"7D",  -- 125
        5285 => X"71",  -- 113
        5286 => X"68",  -- 104
        5287 => X"65",  -- 101
        5288 => X"5B",  -- 91
        5289 => X"59",  -- 89
        5290 => X"56",  -- 86
        5291 => X"58",  -- 88
        5292 => X"59",  -- 89
        5293 => X"5D",  -- 93
        5294 => X"66",  -- 102
        5295 => X"6E",  -- 110
        5296 => X"6E",  -- 110
        5297 => X"6D",  -- 109
        5298 => X"6C",  -- 108
        5299 => X"6B",  -- 107
        5300 => X"6D",  -- 109
        5301 => X"73",  -- 115
        5302 => X"7C",  -- 124
        5303 => X"83",  -- 131
        5304 => X"7A",  -- 122
        5305 => X"78",  -- 120
        5306 => X"77",  -- 119
        5307 => X"79",  -- 121
        5308 => X"7E",  -- 126
        5309 => X"81",  -- 129
        5310 => X"7C",  -- 124
        5311 => X"78",  -- 120
        5312 => X"82",  -- 130
        5313 => X"85",  -- 133
        5314 => X"8E",  -- 142
        5315 => X"93",  -- 147
        5316 => X"8E",  -- 142
        5317 => X"86",  -- 134
        5318 => X"87",  -- 135
        5319 => X"8E",  -- 142
        5320 => X"96",  -- 150
        5321 => X"92",  -- 146
        5322 => X"92",  -- 146
        5323 => X"97",  -- 151
        5324 => X"9A",  -- 154
        5325 => X"99",  -- 153
        5326 => X"9C",  -- 156
        5327 => X"A1",  -- 161
        5328 => X"A8",  -- 168
        5329 => X"AC",  -- 172
        5330 => X"AE",  -- 174
        5331 => X"B3",  -- 179
        5332 => X"B5",  -- 181
        5333 => X"B4",  -- 180
        5334 => X"B4",  -- 180
        5335 => X"B3",  -- 179
        5336 => X"B9",  -- 185
        5337 => X"B9",  -- 185
        5338 => X"B8",  -- 184
        5339 => X"B7",  -- 183
        5340 => X"B7",  -- 183
        5341 => X"B3",  -- 179
        5342 => X"A5",  -- 165
        5343 => X"97",  -- 151
        5344 => X"8F",  -- 143
        5345 => X"88",  -- 136
        5346 => X"86",  -- 134
        5347 => X"85",  -- 133
        5348 => X"89",  -- 137
        5349 => X"95",  -- 149
        5350 => X"99",  -- 153
        5351 => X"8F",  -- 143
        5352 => X"92",  -- 146
        5353 => X"98",  -- 152
        5354 => X"9B",  -- 155
        5355 => X"9A",  -- 154
        5356 => X"98",  -- 152
        5357 => X"9C",  -- 156
        5358 => X"A1",  -- 161
        5359 => X"A3",  -- 163
        5360 => X"A6",  -- 166
        5361 => X"A7",  -- 167
        5362 => X"A5",  -- 165
        5363 => X"A2",  -- 162
        5364 => X"A4",  -- 164
        5365 => X"AA",  -- 170
        5366 => X"AD",  -- 173
        5367 => X"AB",  -- 171
        5368 => X"AF",  -- 175
        5369 => X"B1",  -- 177
        5370 => X"B5",  -- 181
        5371 => X"B7",  -- 183
        5372 => X"B8",  -- 184
        5373 => X"B7",  -- 183
        5374 => X"B6",  -- 182
        5375 => X"B5",  -- 181
        5376 => X"B6",  -- 182
        5377 => X"B6",  -- 182
        5378 => X"B6",  -- 182
        5379 => X"B3",  -- 179
        5380 => X"B1",  -- 177
        5381 => X"AF",  -- 175
        5382 => X"AC",  -- 172
        5383 => X"AA",  -- 170
        5384 => X"A7",  -- 167
        5385 => X"A4",  -- 164
        5386 => X"9F",  -- 159
        5387 => X"98",  -- 152
        5388 => X"97",  -- 151
        5389 => X"9C",  -- 156
        5390 => X"9A",  -- 154
        5391 => X"94",  -- 148
        5392 => X"97",  -- 151
        5393 => X"9B",  -- 155
        5394 => X"9F",  -- 159
        5395 => X"A1",  -- 161
        5396 => X"9B",  -- 155
        5397 => X"94",  -- 148
        5398 => X"8C",  -- 140
        5399 => X"88",  -- 136
        5400 => X"88",  -- 136
        5401 => X"86",  -- 134
        5402 => X"7E",  -- 126
        5403 => X"75",  -- 117
        5404 => X"6D",  -- 109
        5405 => X"63",  -- 99
        5406 => X"53",  -- 83
        5407 => X"47",  -- 71
        5408 => X"5C",  -- 92
        5409 => X"62",  -- 98
        5410 => X"60",  -- 96
        5411 => X"55",  -- 85
        5412 => X"55",  -- 85
        5413 => X"69",  -- 105
        5414 => X"81",  -- 129
        5415 => X"91",  -- 145
        5416 => X"93",  -- 147
        5417 => X"AE",  -- 174
        5418 => X"C0",  -- 192
        5419 => X"C1",  -- 193
        5420 => X"C2",  -- 194
        5421 => X"BF",  -- 191
        5422 => X"BC",  -- 188
        5423 => X"BF",  -- 191
        5424 => X"BF",  -- 191
        5425 => X"C2",  -- 194
        5426 => X"C3",  -- 195
        5427 => X"C2",  -- 194
        5428 => X"C0",  -- 192
        5429 => X"BC",  -- 188
        5430 => X"B7",  -- 183
        5431 => X"B4",  -- 180
        5432 => X"B2",  -- 178
        5433 => X"AF",  -- 175
        5434 => X"B1",  -- 177
        5435 => X"B8",  -- 184
        5436 => X"B7",  -- 183
        5437 => X"B3",  -- 179
        5438 => X"B7",  -- 183
        5439 => X"C0",  -- 192
        5440 => X"3F",  -- 63
        5441 => X"3E",  -- 62
        5442 => X"3D",  -- 61
        5443 => X"3B",  -- 59
        5444 => X"3A",  -- 58
        5445 => X"3A",  -- 58
        5446 => X"3A",  -- 58
        5447 => X"3A",  -- 58
        5448 => X"3A",  -- 58
        5449 => X"3A",  -- 58
        5450 => X"3B",  -- 59
        5451 => X"3B",  -- 59
        5452 => X"3C",  -- 60
        5453 => X"3C",  -- 60
        5454 => X"3D",  -- 61
        5455 => X"3D",  -- 61
        5456 => X"3D",  -- 61
        5457 => X"3D",  -- 61
        5458 => X"3D",  -- 61
        5459 => X"3D",  -- 61
        5460 => X"3D",  -- 61
        5461 => X"3D",  -- 61
        5462 => X"3D",  -- 61
        5463 => X"3D",  -- 61
        5464 => X"3D",  -- 61
        5465 => X"3E",  -- 62
        5466 => X"3F",  -- 63
        5467 => X"40",  -- 64
        5468 => X"40",  -- 64
        5469 => X"41",  -- 65
        5470 => X"40",  -- 64
        5471 => X"40",  -- 64
        5472 => X"3E",  -- 62
        5473 => X"3E",  -- 62
        5474 => X"3D",  -- 61
        5475 => X"3B",  -- 59
        5476 => X"3B",  -- 59
        5477 => X"3A",  -- 58
        5478 => X"39",  -- 57
        5479 => X"38",  -- 56
        5480 => X"36",  -- 54
        5481 => X"35",  -- 53
        5482 => X"35",  -- 53
        5483 => X"34",  -- 52
        5484 => X"33",  -- 51
        5485 => X"33",  -- 51
        5486 => X"32",  -- 50
        5487 => X"32",  -- 50
        5488 => X"31",  -- 49
        5489 => X"31",  -- 49
        5490 => X"31",  -- 49
        5491 => X"30",  -- 48
        5492 => X"2E",  -- 46
        5493 => X"2E",  -- 46
        5494 => X"2D",  -- 45
        5495 => X"2D",  -- 45
        5496 => X"2F",  -- 47
        5497 => X"2D",  -- 45
        5498 => X"2C",  -- 44
        5499 => X"2A",  -- 42
        5500 => X"2B",  -- 43
        5501 => X"2B",  -- 43
        5502 => X"29",  -- 41
        5503 => X"28",  -- 40
        5504 => X"2B",  -- 43
        5505 => X"2E",  -- 46
        5506 => X"32",  -- 50
        5507 => X"36",  -- 54
        5508 => X"3A",  -- 58
        5509 => X"3D",  -- 61
        5510 => X"40",  -- 64
        5511 => X"41",  -- 65
        5512 => X"43",  -- 67
        5513 => X"45",  -- 69
        5514 => X"47",  -- 71
        5515 => X"47",  -- 71
        5516 => X"48",  -- 72
        5517 => X"4B",  -- 75
        5518 => X"51",  -- 81
        5519 => X"56",  -- 86
        5520 => X"5D",  -- 93
        5521 => X"6A",  -- 106
        5522 => X"79",  -- 121
        5523 => X"94",  -- 148
        5524 => X"A1",  -- 161
        5525 => X"9D",  -- 157
        5526 => X"A4",  -- 164
        5527 => X"A5",  -- 165
        5528 => X"A3",  -- 163
        5529 => X"A6",  -- 166
        5530 => X"A3",  -- 163
        5531 => X"9A",  -- 154
        5532 => X"9A",  -- 154
        5533 => X"A3",  -- 163
        5534 => X"A7",  -- 167
        5535 => X"A2",  -- 162
        5536 => X"9C",  -- 156
        5537 => X"98",  -- 152
        5538 => X"9D",  -- 157
        5539 => X"96",  -- 150
        5540 => X"94",  -- 148
        5541 => X"98",  -- 152
        5542 => X"8E",  -- 142
        5543 => X"90",  -- 144
        5544 => X"86",  -- 134
        5545 => X"7A",  -- 122
        5546 => X"6E",  -- 110
        5547 => X"53",  -- 83
        5548 => X"46",  -- 70
        5549 => X"35",  -- 53
        5550 => X"41",  -- 65
        5551 => X"4A",  -- 74
        5552 => X"68",  -- 104
        5553 => X"6E",  -- 110
        5554 => X"6F",  -- 111
        5555 => X"78",  -- 120
        5556 => X"6E",  -- 110
        5557 => X"83",  -- 131
        5558 => X"8A",  -- 138
        5559 => X"8B",  -- 139
        5560 => X"90",  -- 144
        5561 => X"8E",  -- 142
        5562 => X"8E",  -- 142
        5563 => X"91",  -- 145
        5564 => X"93",  -- 147
        5565 => X"93",  -- 147
        5566 => X"8F",  -- 143
        5567 => X"8B",  -- 139
        5568 => X"8C",  -- 140
        5569 => X"90",  -- 144
        5570 => X"8D",  -- 141
        5571 => X"7B",  -- 123
        5572 => X"68",  -- 104
        5573 => X"67",  -- 103
        5574 => X"65",  -- 101
        5575 => X"5B",  -- 91
        5576 => X"6A",  -- 106
        5577 => X"58",  -- 88
        5578 => X"4B",  -- 75
        5579 => X"4D",  -- 77
        5580 => X"49",  -- 73
        5581 => X"36",  -- 54
        5582 => X"37",  -- 55
        5583 => X"4E",  -- 78
        5584 => X"4B",  -- 75
        5585 => X"46",  -- 70
        5586 => X"45",  -- 69
        5587 => X"4A",  -- 74
        5588 => X"58",  -- 88
        5589 => X"5E",  -- 94
        5590 => X"58",  -- 88
        5591 => X"50",  -- 80
        5592 => X"4E",  -- 78
        5593 => X"4C",  -- 76
        5594 => X"45",  -- 69
        5595 => X"40",  -- 64
        5596 => X"43",  -- 67
        5597 => X"50",  -- 80
        5598 => X"5C",  -- 92
        5599 => X"62",  -- 98
        5600 => X"7C",  -- 124
        5601 => X"88",  -- 136
        5602 => X"92",  -- 146
        5603 => X"90",  -- 144
        5604 => X"87",  -- 135
        5605 => X"7E",  -- 126
        5606 => X"7A",  -- 122
        5607 => X"75",  -- 117
        5608 => X"5F",  -- 95
        5609 => X"56",  -- 86
        5610 => X"4E",  -- 78
        5611 => X"51",  -- 81
        5612 => X"58",  -- 88
        5613 => X"5C",  -- 92
        5614 => X"60",  -- 96
        5615 => X"63",  -- 99
        5616 => X"62",  -- 98
        5617 => X"67",  -- 103
        5618 => X"6D",  -- 109
        5619 => X"70",  -- 112
        5620 => X"72",  -- 114
        5621 => X"71",  -- 113
        5622 => X"70",  -- 112
        5623 => X"71",  -- 113
        5624 => X"74",  -- 116
        5625 => X"74",  -- 116
        5626 => X"75",  -- 117
        5627 => X"76",  -- 118
        5628 => X"79",  -- 121
        5629 => X"7C",  -- 124
        5630 => X"80",  -- 128
        5631 => X"81",  -- 129
        5632 => X"7D",  -- 125
        5633 => X"80",  -- 128
        5634 => X"89",  -- 137
        5635 => X"90",  -- 144
        5636 => X"90",  -- 144
        5637 => X"8E",  -- 142
        5638 => X"90",  -- 144
        5639 => X"97",  -- 151
        5640 => X"91",  -- 145
        5641 => X"92",  -- 146
        5642 => X"96",  -- 150
        5643 => X"9A",  -- 154
        5644 => X"99",  -- 153
        5645 => X"98",  -- 152
        5646 => X"9D",  -- 157
        5647 => X"A4",  -- 164
        5648 => X"A6",  -- 166
        5649 => X"A9",  -- 169
        5650 => X"AC",  -- 172
        5651 => X"AF",  -- 175
        5652 => X"B3",  -- 179
        5653 => X"B5",  -- 181
        5654 => X"B6",  -- 182
        5655 => X"B6",  -- 182
        5656 => X"B8",  -- 184
        5657 => X"B7",  -- 183
        5658 => X"B6",  -- 182
        5659 => X"B5",  -- 181
        5660 => X"B5",  -- 181
        5661 => X"B1",  -- 177
        5662 => X"A5",  -- 165
        5663 => X"97",  -- 151
        5664 => X"8E",  -- 142
        5665 => X"83",  -- 131
        5666 => X"80",  -- 128
        5667 => X"83",  -- 131
        5668 => X"86",  -- 134
        5669 => X"8C",  -- 140
        5670 => X"8D",  -- 141
        5671 => X"86",  -- 134
        5672 => X"90",  -- 144
        5673 => X"97",  -- 151
        5674 => X"9C",  -- 156
        5675 => X"9B",  -- 155
        5676 => X"9B",  -- 155
        5677 => X"9E",  -- 158
        5678 => X"A4",  -- 164
        5679 => X"A5",  -- 165
        5680 => X"AC",  -- 172
        5681 => X"AD",  -- 173
        5682 => X"AC",  -- 172
        5683 => X"A9",  -- 169
        5684 => X"AA",  -- 170
        5685 => X"AD",  -- 173
        5686 => X"AE",  -- 174
        5687 => X"AB",  -- 171
        5688 => X"AD",  -- 173
        5689 => X"B0",  -- 176
        5690 => X"B5",  -- 181
        5691 => X"B9",  -- 185
        5692 => X"BA",  -- 186
        5693 => X"B9",  -- 185
        5694 => X"B7",  -- 183
        5695 => X"B5",  -- 181
        5696 => X"B5",  -- 181
        5697 => X"B6",  -- 182
        5698 => X"B4",  -- 180
        5699 => X"B4",  -- 180
        5700 => X"B4",  -- 180
        5701 => X"B0",  -- 176
        5702 => X"AA",  -- 170
        5703 => X"A8",  -- 168
        5704 => X"9E",  -- 158
        5705 => X"9C",  -- 156
        5706 => X"9E",  -- 158
        5707 => X"9C",  -- 156
        5708 => X"95",  -- 149
        5709 => X"99",  -- 153
        5710 => X"9D",  -- 157
        5711 => X"97",  -- 151
        5712 => X"96",  -- 150
        5713 => X"98",  -- 152
        5714 => X"9B",  -- 155
        5715 => X"9E",  -- 158
        5716 => X"9C",  -- 156
        5717 => X"9A",  -- 154
        5718 => X"98",  -- 152
        5719 => X"96",  -- 150
        5720 => X"95",  -- 149
        5721 => X"91",  -- 145
        5722 => X"87",  -- 135
        5723 => X"7B",  -- 123
        5724 => X"73",  -- 115
        5725 => X"6C",  -- 108
        5726 => X"61",  -- 97
        5727 => X"57",  -- 87
        5728 => X"5E",  -- 94
        5729 => X"58",  -- 88
        5730 => X"4E",  -- 78
        5731 => X"4B",  -- 75
        5732 => X"57",  -- 87
        5733 => X"6B",  -- 107
        5734 => X"77",  -- 119
        5735 => X"7B",  -- 123
        5736 => X"8A",  -- 138
        5737 => X"A6",  -- 166
        5738 => X"BA",  -- 186
        5739 => X"BE",  -- 190
        5740 => X"C1",  -- 193
        5741 => X"C1",  -- 193
        5742 => X"BE",  -- 190
        5743 => X"C0",  -- 192
        5744 => X"BE",  -- 190
        5745 => X"BF",  -- 191
        5746 => X"BF",  -- 191
        5747 => X"C0",  -- 192
        5748 => X"BF",  -- 191
        5749 => X"BF",  -- 191
        5750 => X"C0",  -- 192
        5751 => X"C0",  -- 192
        5752 => X"B8",  -- 184
        5753 => X"B4",  -- 180
        5754 => X"B3",  -- 179
        5755 => X"B5",  -- 181
        5756 => X"B3",  -- 179
        5757 => X"AF",  -- 175
        5758 => X"B4",  -- 180
        5759 => X"BF",  -- 191
        5760 => X"3E",  -- 62
        5761 => X"3E",  -- 62
        5762 => X"3C",  -- 60
        5763 => X"3B",  -- 59
        5764 => X"3A",  -- 58
        5765 => X"3A",  -- 58
        5766 => X"3A",  -- 58
        5767 => X"3A",  -- 58
        5768 => X"3A",  -- 58
        5769 => X"3B",  -- 59
        5770 => X"3B",  -- 59
        5771 => X"3B",  -- 59
        5772 => X"3C",  -- 60
        5773 => X"3D",  -- 61
        5774 => X"3D",  -- 61
        5775 => X"3D",  -- 61
        5776 => X"3D",  -- 61
        5777 => X"3D",  -- 61
        5778 => X"3D",  -- 61
        5779 => X"3D",  -- 61
        5780 => X"3D",  -- 61
        5781 => X"3D",  -- 61
        5782 => X"3D",  -- 61
        5783 => X"3D",  -- 61
        5784 => X"3D",  -- 61
        5785 => X"3E",  -- 62
        5786 => X"3E",  -- 62
        5787 => X"3F",  -- 63
        5788 => X"40",  -- 64
        5789 => X"40",  -- 64
        5790 => X"40",  -- 64
        5791 => X"40",  -- 64
        5792 => X"3E",  -- 62
        5793 => X"3D",  -- 61
        5794 => X"3C",  -- 60
        5795 => X"3B",  -- 59
        5796 => X"3A",  -- 58
        5797 => X"39",  -- 57
        5798 => X"39",  -- 57
        5799 => X"38",  -- 56
        5800 => X"36",  -- 54
        5801 => X"36",  -- 54
        5802 => X"34",  -- 52
        5803 => X"34",  -- 52
        5804 => X"33",  -- 51
        5805 => X"32",  -- 50
        5806 => X"31",  -- 49
        5807 => X"31",  -- 49
        5808 => X"32",  -- 50
        5809 => X"32",  -- 50
        5810 => X"31",  -- 49
        5811 => X"2F",  -- 47
        5812 => X"2F",  -- 47
        5813 => X"2E",  -- 46
        5814 => X"2D",  -- 45
        5815 => X"2D",  -- 45
        5816 => X"2C",  -- 44
        5817 => X"2C",  -- 44
        5818 => X"2B",  -- 43
        5819 => X"2A",  -- 42
        5820 => X"2A",  -- 42
        5821 => X"2A",  -- 42
        5822 => X"28",  -- 40
        5823 => X"28",  -- 40
        5824 => X"2A",  -- 42
        5825 => X"2E",  -- 46
        5826 => X"32",  -- 50
        5827 => X"35",  -- 53
        5828 => X"38",  -- 56
        5829 => X"3A",  -- 58
        5830 => X"3D",  -- 61
        5831 => X"3F",  -- 63
        5832 => X"43",  -- 67
        5833 => X"46",  -- 70
        5834 => X"4A",  -- 74
        5835 => X"4C",  -- 76
        5836 => X"4E",  -- 78
        5837 => X"53",  -- 83
        5838 => X"5D",  -- 93
        5839 => X"65",  -- 101
        5840 => X"76",  -- 118
        5841 => X"84",  -- 132
        5842 => X"8D",  -- 141
        5843 => X"9F",  -- 159
        5844 => X"A9",  -- 169
        5845 => X"A5",  -- 165
        5846 => X"A5",  -- 165
        5847 => X"9C",  -- 156
        5848 => X"9B",  -- 155
        5849 => X"A5",  -- 165
        5850 => X"A5",  -- 165
        5851 => X"9A",  -- 154
        5852 => X"98",  -- 152
        5853 => X"A1",  -- 161
        5854 => X"A3",  -- 163
        5855 => X"9D",  -- 157
        5856 => X"9D",  -- 157
        5857 => X"9E",  -- 158
        5858 => X"A0",  -- 160
        5859 => X"93",  -- 147
        5860 => X"8F",  -- 143
        5861 => X"99",  -- 153
        5862 => X"92",  -- 146
        5863 => X"8F",  -- 143
        5864 => X"86",  -- 134
        5865 => X"76",  -- 118
        5866 => X"6D",  -- 109
        5867 => X"55",  -- 85
        5868 => X"46",  -- 70
        5869 => X"31",  -- 49
        5870 => X"41",  -- 65
        5871 => X"51",  -- 81
        5872 => X"62",  -- 98
        5873 => X"62",  -- 98
        5874 => X"5C",  -- 92
        5875 => X"5D",  -- 93
        5876 => X"5E",  -- 94
        5877 => X"7F",  -- 127
        5878 => X"8C",  -- 140
        5879 => X"87",  -- 135
        5880 => X"89",  -- 137
        5881 => X"8C",  -- 140
        5882 => X"8F",  -- 143
        5883 => X"92",  -- 146
        5884 => X"91",  -- 145
        5885 => X"90",  -- 144
        5886 => X"8D",  -- 141
        5887 => X"8A",  -- 138
        5888 => X"90",  -- 144
        5889 => X"93",  -- 147
        5890 => X"88",  -- 136
        5891 => X"78",  -- 120
        5892 => X"71",  -- 113
        5893 => X"68",  -- 104
        5894 => X"62",  -- 98
        5895 => X"62",  -- 98
        5896 => X"67",  -- 103
        5897 => X"4B",  -- 75
        5898 => X"41",  -- 65
        5899 => X"4C",  -- 76
        5900 => X"43",  -- 67
        5901 => X"36",  -- 54
        5902 => X"3F",  -- 63
        5903 => X"53",  -- 83
        5904 => X"53",  -- 83
        5905 => X"4A",  -- 74
        5906 => X"4C",  -- 76
        5907 => X"58",  -- 88
        5908 => X"5E",  -- 94
        5909 => X"54",  -- 84
        5910 => X"4D",  -- 77
        5911 => X"51",  -- 81
        5912 => X"51",  -- 81
        5913 => X"59",  -- 89
        5914 => X"5E",  -- 94
        5915 => X"5B",  -- 91
        5916 => X"57",  -- 87
        5917 => X"56",  -- 86
        5918 => X"57",  -- 87
        5919 => X"56",  -- 86
        5920 => X"5F",  -- 95
        5921 => X"6A",  -- 106
        5922 => X"77",  -- 119
        5923 => X"7E",  -- 126
        5924 => X"7D",  -- 125
        5925 => X"7A",  -- 122
        5926 => X"72",  -- 114
        5927 => X"6D",  -- 109
        5928 => X"56",  -- 86
        5929 => X"49",  -- 73
        5930 => X"40",  -- 64
        5931 => X"47",  -- 71
        5932 => X"56",  -- 86
        5933 => X"5F",  -- 95
        5934 => X"61",  -- 97
        5935 => X"5F",  -- 95
        5936 => X"62",  -- 98
        5937 => X"68",  -- 104
        5938 => X"70",  -- 112
        5939 => X"74",  -- 116
        5940 => X"76",  -- 118
        5941 => X"72",  -- 114
        5942 => X"6D",  -- 109
        5943 => X"6B",  -- 107
        5944 => X"78",  -- 120
        5945 => X"78",  -- 120
        5946 => X"75",  -- 117
        5947 => X"73",  -- 115
        5948 => X"72",  -- 114
        5949 => X"75",  -- 117
        5950 => X"7D",  -- 125
        5951 => X"81",  -- 129
        5952 => X"85",  -- 133
        5953 => X"86",  -- 134
        5954 => X"88",  -- 136
        5955 => X"8B",  -- 139
        5956 => X"8C",  -- 140
        5957 => X"8B",  -- 139
        5958 => X"8B",  -- 139
        5959 => X"8F",  -- 143
        5960 => X"8E",  -- 142
        5961 => X"93",  -- 147
        5962 => X"9A",  -- 154
        5963 => X"9C",  -- 156
        5964 => X"98",  -- 152
        5965 => X"97",  -- 151
        5966 => X"9C",  -- 156
        5967 => X"A4",  -- 164
        5968 => X"A4",  -- 164
        5969 => X"A6",  -- 166
        5970 => X"A9",  -- 169
        5971 => X"AD",  -- 173
        5972 => X"B0",  -- 176
        5973 => X"B3",  -- 179
        5974 => X"B6",  -- 182
        5975 => X"B8",  -- 184
        5976 => X"B9",  -- 185
        5977 => X"B8",  -- 184
        5978 => X"B6",  -- 182
        5979 => X"B4",  -- 180
        5980 => X"B4",  -- 180
        5981 => X"B1",  -- 177
        5982 => X"A7",  -- 167
        5983 => X"9B",  -- 155
        5984 => X"8D",  -- 141
        5985 => X"7F",  -- 127
        5986 => X"7F",  -- 127
        5987 => X"87",  -- 135
        5988 => X"8A",  -- 138
        5989 => X"8A",  -- 138
        5990 => X"8B",  -- 139
        5991 => X"89",  -- 137
        5992 => X"8F",  -- 143
        5993 => X"96",  -- 150
        5994 => X"9B",  -- 155
        5995 => X"9C",  -- 156
        5996 => X"9D",  -- 157
        5997 => X"A1",  -- 161
        5998 => X"A5",  -- 165
        5999 => X"A6",  -- 166
        6000 => X"A7",  -- 167
        6001 => X"AB",  -- 171
        6002 => X"AC",  -- 172
        6003 => X"AB",  -- 171
        6004 => X"AB",  -- 171
        6005 => X"AB",  -- 171
        6006 => X"A9",  -- 169
        6007 => X"A6",  -- 166
        6008 => X"AA",  -- 170
        6009 => X"AE",  -- 174
        6010 => X"B3",  -- 179
        6011 => X"B8",  -- 184
        6012 => X"BB",  -- 187
        6013 => X"BA",  -- 186
        6014 => X"B7",  -- 183
        6015 => X"B5",  -- 181
        6016 => X"B4",  -- 180
        6017 => X"B3",  -- 179
        6018 => X"B3",  -- 179
        6019 => X"B5",  -- 181
        6020 => X"B7",  -- 183
        6021 => X"B1",  -- 177
        6022 => X"A8",  -- 168
        6023 => X"A2",  -- 162
        6024 => X"95",  -- 149
        6025 => X"91",  -- 145
        6026 => X"9B",  -- 155
        6027 => X"9D",  -- 157
        6028 => X"91",  -- 145
        6029 => X"97",  -- 151
        6030 => X"9E",  -- 158
        6031 => X"96",  -- 150
        6032 => X"9C",  -- 156
        6033 => X"9D",  -- 157
        6034 => X"9C",  -- 156
        6035 => X"9A",  -- 154
        6036 => X"98",  -- 152
        6037 => X"97",  -- 151
        6038 => X"99",  -- 153
        6039 => X"9A",  -- 154
        6040 => X"99",  -- 153
        6041 => X"96",  -- 150
        6042 => X"8E",  -- 142
        6043 => X"84",  -- 132
        6044 => X"7B",  -- 123
        6045 => X"74",  -- 116
        6046 => X"66",  -- 102
        6047 => X"5B",  -- 91
        6048 => X"53",  -- 83
        6049 => X"4D",  -- 77
        6050 => X"47",  -- 71
        6051 => X"4A",  -- 74
        6052 => X"58",  -- 88
        6053 => X"65",  -- 101
        6054 => X"69",  -- 105
        6055 => X"67",  -- 103
        6056 => X"85",  -- 133
        6057 => X"A1",  -- 161
        6058 => X"B4",  -- 180
        6059 => X"B8",  -- 184
        6060 => X"BB",  -- 187
        6061 => X"BC",  -- 188
        6062 => X"B9",  -- 185
        6063 => X"BB",  -- 187
        6064 => X"BB",  -- 187
        6065 => X"BA",  -- 186
        6066 => X"BB",  -- 187
        6067 => X"BB",  -- 187
        6068 => X"BC",  -- 188
        6069 => X"BF",  -- 191
        6070 => X"C1",  -- 193
        6071 => X"C4",  -- 196
        6072 => X"BF",  -- 191
        6073 => X"BA",  -- 186
        6074 => X"B6",  -- 182
        6075 => X"B4",  -- 180
        6076 => X"AE",  -- 174
        6077 => X"A9",  -- 169
        6078 => X"AD",  -- 173
        6079 => X"B9",  -- 185
        6080 => X"3E",  -- 62
        6081 => X"3D",  -- 61
        6082 => X"3C",  -- 60
        6083 => X"3B",  -- 59
        6084 => X"3B",  -- 59
        6085 => X"3A",  -- 58
        6086 => X"3A",  -- 58
        6087 => X"3B",  -- 59
        6088 => X"3B",  -- 59
        6089 => X"3B",  -- 59
        6090 => X"3B",  -- 59
        6091 => X"3C",  -- 60
        6092 => X"3C",  -- 60
        6093 => X"3D",  -- 61
        6094 => X"3D",  -- 61
        6095 => X"3D",  -- 61
        6096 => X"3D",  -- 61
        6097 => X"3D",  -- 61
        6098 => X"3D",  -- 61
        6099 => X"3D",  -- 61
        6100 => X"3D",  -- 61
        6101 => X"3D",  -- 61
        6102 => X"3D",  -- 61
        6103 => X"3D",  -- 61
        6104 => X"3D",  -- 61
        6105 => X"3E",  -- 62
        6106 => X"3E",  -- 62
        6107 => X"3F",  -- 63
        6108 => X"40",  -- 64
        6109 => X"3F",  -- 63
        6110 => X"3F",  -- 63
        6111 => X"3F",  -- 63
        6112 => X"3E",  -- 62
        6113 => X"3D",  -- 61
        6114 => X"3C",  -- 60
        6115 => X"3B",  -- 59
        6116 => X"39",  -- 57
        6117 => X"38",  -- 56
        6118 => X"38",  -- 56
        6119 => X"38",  -- 56
        6120 => X"36",  -- 54
        6121 => X"36",  -- 54
        6122 => X"34",  -- 52
        6123 => X"34",  -- 52
        6124 => X"34",  -- 52
        6125 => X"32",  -- 50
        6126 => X"33",  -- 51
        6127 => X"32",  -- 50
        6128 => X"31",  -- 49
        6129 => X"31",  -- 49
        6130 => X"30",  -- 48
        6131 => X"30",  -- 48
        6132 => X"30",  -- 48
        6133 => X"2E",  -- 46
        6134 => X"2F",  -- 47
        6135 => X"2D",  -- 45
        6136 => X"29",  -- 41
        6137 => X"2A",  -- 42
        6138 => X"2A",  -- 42
        6139 => X"2A",  -- 42
        6140 => X"2B",  -- 43
        6141 => X"2A",  -- 42
        6142 => X"2A",  -- 42
        6143 => X"2A",  -- 42
        6144 => X"2D",  -- 45
        6145 => X"2F",  -- 47
        6146 => X"32",  -- 50
        6147 => X"33",  -- 51
        6148 => X"37",  -- 55
        6149 => X"3A",  -- 58
        6150 => X"3E",  -- 62
        6151 => X"42",  -- 66
        6152 => X"48",  -- 72
        6153 => X"4D",  -- 77
        6154 => X"54",  -- 84
        6155 => X"59",  -- 89
        6156 => X"5B",  -- 91
        6157 => X"63",  -- 99
        6158 => X"6F",  -- 111
        6159 => X"76",  -- 118
        6160 => X"8E",  -- 142
        6161 => X"9C",  -- 156
        6162 => X"9D",  -- 157
        6163 => X"A4",  -- 164
        6164 => X"A7",  -- 167
        6165 => X"A2",  -- 162
        6166 => X"A6",  -- 166
        6167 => X"9C",  -- 156
        6168 => X"96",  -- 150
        6169 => X"A3",  -- 163
        6170 => X"A5",  -- 165
        6171 => X"9B",  -- 155
        6172 => X"98",  -- 152
        6173 => X"A0",  -- 160
        6174 => X"A2",  -- 162
        6175 => X"9D",  -- 157
        6176 => X"9B",  -- 155
        6177 => X"9B",  -- 155
        6178 => X"A4",  -- 164
        6179 => X"9A",  -- 154
        6180 => X"97",  -- 151
        6181 => X"9B",  -- 155
        6182 => X"8F",  -- 143
        6183 => X"8C",  -- 140
        6184 => X"82",  -- 130
        6185 => X"77",  -- 119
        6186 => X"74",  -- 116
        6187 => X"60",  -- 96
        6188 => X"4F",  -- 79
        6189 => X"34",  -- 52
        6190 => X"42",  -- 66
        6191 => X"55",  -- 85
        6192 => X"56",  -- 86
        6193 => X"4C",  -- 76
        6194 => X"45",  -- 69
        6195 => X"49",  -- 73
        6196 => X"54",  -- 84
        6197 => X"74",  -- 116
        6198 => X"86",  -- 134
        6199 => X"87",  -- 135
        6200 => X"84",  -- 132
        6201 => X"88",  -- 136
        6202 => X"8E",  -- 142
        6203 => X"90",  -- 144
        6204 => X"90",  -- 144
        6205 => X"8F",  -- 143
        6206 => X"8F",  -- 143
        6207 => X"8F",  -- 143
        6208 => X"8D",  -- 141
        6209 => X"90",  -- 144
        6210 => X"86",  -- 134
        6211 => X"80",  -- 128
        6212 => X"7F",  -- 127
        6213 => X"6C",  -- 108
        6214 => X"58",  -- 88
        6215 => X"59",  -- 89
        6216 => X"52",  -- 82
        6217 => X"39",  -- 57
        6218 => X"39",  -- 57
        6219 => X"46",  -- 70
        6220 => X"3F",  -- 63
        6221 => X"3C",  -- 60
        6222 => X"4A",  -- 74
        6223 => X"55",  -- 85
        6224 => X"4D",  -- 77
        6225 => X"4B",  -- 75
        6226 => X"53",  -- 83
        6227 => X"5E",  -- 94
        6228 => X"57",  -- 87
        6229 => X"46",  -- 70
        6230 => X"40",  -- 64
        6231 => X"46",  -- 70
        6232 => X"4A",  -- 74
        6233 => X"55",  -- 85
        6234 => X"5F",  -- 95
        6235 => X"61",  -- 97
        6236 => X"60",  -- 96
        6237 => X"5E",  -- 94
        6238 => X"58",  -- 88
        6239 => X"51",  -- 81
        6240 => X"55",  -- 85
        6241 => X"5C",  -- 92
        6242 => X"6A",  -- 106
        6243 => X"77",  -- 119
        6244 => X"7E",  -- 126
        6245 => X"7A",  -- 122
        6246 => X"6D",  -- 109
        6247 => X"61",  -- 97
        6248 => X"45",  -- 69
        6249 => X"3C",  -- 60
        6250 => X"38",  -- 56
        6251 => X"42",  -- 66
        6252 => X"55",  -- 85
        6253 => X"62",  -- 98
        6254 => X"66",  -- 102
        6255 => X"64",  -- 100
        6256 => X"6B",  -- 107
        6257 => X"6C",  -- 108
        6258 => X"6D",  -- 109
        6259 => X"6F",  -- 111
        6260 => X"70",  -- 112
        6261 => X"71",  -- 113
        6262 => X"71",  -- 113
        6263 => X"71",  -- 113
        6264 => X"77",  -- 119
        6265 => X"75",  -- 117
        6266 => X"73",  -- 115
        6267 => X"72",  -- 114
        6268 => X"73",  -- 115
        6269 => X"77",  -- 119
        6270 => X"7D",  -- 125
        6271 => X"80",  -- 128
        6272 => X"8B",  -- 139
        6273 => X"88",  -- 136
        6274 => X"86",  -- 134
        6275 => X"85",  -- 133
        6276 => X"85",  -- 133
        6277 => X"85",  -- 133
        6278 => X"84",  -- 132
        6279 => X"84",  -- 132
        6280 => X"91",  -- 145
        6281 => X"94",  -- 148
        6282 => X"98",  -- 152
        6283 => X"98",  -- 152
        6284 => X"95",  -- 149
        6285 => X"95",  -- 149
        6286 => X"9B",  -- 155
        6287 => X"A1",  -- 161
        6288 => X"A4",  -- 164
        6289 => X"A5",  -- 165
        6290 => X"A8",  -- 168
        6291 => X"AB",  -- 171
        6292 => X"AE",  -- 174
        6293 => X"B2",  -- 178
        6294 => X"B6",  -- 182
        6295 => X"B8",  -- 184
        6296 => X"BB",  -- 187
        6297 => X"BA",  -- 186
        6298 => X"B9",  -- 185
        6299 => X"B6",  -- 182
        6300 => X"B5",  -- 181
        6301 => X"B4",  -- 180
        6302 => X"AC",  -- 172
        6303 => X"A2",  -- 162
        6304 => X"8B",  -- 139
        6305 => X"7C",  -- 124
        6306 => X"7D",  -- 125
        6307 => X"8C",  -- 140
        6308 => X"8F",  -- 143
        6309 => X"8C",  -- 140
        6310 => X"8F",  -- 143
        6311 => X"91",  -- 145
        6312 => X"8F",  -- 143
        6313 => X"96",  -- 150
        6314 => X"99",  -- 153
        6315 => X"9B",  -- 155
        6316 => X"9B",  -- 155
        6317 => X"A0",  -- 160
        6318 => X"A4",  -- 164
        6319 => X"A3",  -- 163
        6320 => X"9F",  -- 159
        6321 => X"A5",  -- 165
        6322 => X"AA",  -- 170
        6323 => X"AB",  -- 171
        6324 => X"AB",  -- 171
        6325 => X"AB",  -- 171
        6326 => X"A8",  -- 168
        6327 => X"A4",  -- 164
        6328 => X"AB",  -- 171
        6329 => X"AD",  -- 173
        6330 => X"B1",  -- 177
        6331 => X"B4",  -- 180
        6332 => X"B7",  -- 183
        6333 => X"B7",  -- 183
        6334 => X"B5",  -- 181
        6335 => X"B3",  -- 179
        6336 => X"B5",  -- 181
        6337 => X"B3",  -- 179
        6338 => X"B3",  -- 179
        6339 => X"B5",  -- 181
        6340 => X"B7",  -- 183
        6341 => X"B1",  -- 177
        6342 => X"A5",  -- 165
        6343 => X"9A",  -- 154
        6344 => X"90",  -- 144
        6345 => X"87",  -- 135
        6346 => X"90",  -- 144
        6347 => X"95",  -- 149
        6348 => X"8D",  -- 141
        6349 => X"94",  -- 148
        6350 => X"A0",  -- 160
        6351 => X"97",  -- 151
        6352 => X"9D",  -- 157
        6353 => X"9E",  -- 158
        6354 => X"9C",  -- 156
        6355 => X"99",  -- 153
        6356 => X"97",  -- 151
        6357 => X"96",  -- 150
        6358 => X"96",  -- 150
        6359 => X"98",  -- 152
        6360 => X"96",  -- 150
        6361 => X"96",  -- 150
        6362 => X"94",  -- 148
        6363 => X"8F",  -- 143
        6364 => X"88",  -- 136
        6365 => X"7D",  -- 125
        6366 => X"6B",  -- 107
        6367 => X"5D",  -- 93
        6368 => X"4F",  -- 79
        6369 => X"50",  -- 80
        6370 => X"53",  -- 83
        6371 => X"56",  -- 86
        6372 => X"56",  -- 86
        6373 => X"54",  -- 84
        6374 => X"54",  -- 84
        6375 => X"56",  -- 86
        6376 => X"7C",  -- 124
        6377 => X"98",  -- 152
        6378 => X"AC",  -- 172
        6379 => X"B3",  -- 179
        6380 => X"B8",  -- 184
        6381 => X"BA",  -- 186
        6382 => X"B7",  -- 183
        6383 => X"BA",  -- 186
        6384 => X"BC",  -- 188
        6385 => X"BB",  -- 187
        6386 => X"B9",  -- 185
        6387 => X"B8",  -- 184
        6388 => X"B9",  -- 185
        6389 => X"BB",  -- 187
        6390 => X"BD",  -- 189
        6391 => X"BF",  -- 191
        6392 => X"C3",  -- 195
        6393 => X"BF",  -- 191
        6394 => X"BA",  -- 186
        6395 => X"B3",  -- 179
        6396 => X"AA",  -- 170
        6397 => X"A3",  -- 163
        6398 => X"A8",  -- 168
        6399 => X"AF",  -- 175
        6400 => X"3D",  -- 61
        6401 => X"3D",  -- 61
        6402 => X"3C",  -- 60
        6403 => X"3B",  -- 59
        6404 => X"3B",  -- 59
        6405 => X"3B",  -- 59
        6406 => X"3B",  -- 59
        6407 => X"3B",  -- 59
        6408 => X"3B",  -- 59
        6409 => X"3B",  -- 59
        6410 => X"3C",  -- 60
        6411 => X"3C",  -- 60
        6412 => X"3D",  -- 61
        6413 => X"3D",  -- 61
        6414 => X"3E",  -- 62
        6415 => X"3E",  -- 62
        6416 => X"3D",  -- 61
        6417 => X"3D",  -- 61
        6418 => X"3D",  -- 61
        6419 => X"3D",  -- 61
        6420 => X"3D",  -- 61
        6421 => X"3D",  -- 61
        6422 => X"3D",  -- 61
        6423 => X"3D",  -- 61
        6424 => X"3D",  -- 61
        6425 => X"3E",  -- 62
        6426 => X"3E",  -- 62
        6427 => X"3F",  -- 63
        6428 => X"3F",  -- 63
        6429 => X"3F",  -- 63
        6430 => X"3E",  -- 62
        6431 => X"3E",  -- 62
        6432 => X"3E",  -- 62
        6433 => X"3D",  -- 61
        6434 => X"3D",  -- 61
        6435 => X"3C",  -- 60
        6436 => X"3A",  -- 58
        6437 => X"39",  -- 57
        6438 => X"38",  -- 56
        6439 => X"37",  -- 55
        6440 => X"34",  -- 52
        6441 => X"34",  -- 52
        6442 => X"34",  -- 52
        6443 => X"33",  -- 51
        6444 => X"33",  -- 51
        6445 => X"33",  -- 51
        6446 => X"32",  -- 50
        6447 => X"32",  -- 50
        6448 => X"33",  -- 51
        6449 => X"32",  -- 50
        6450 => X"32",  -- 50
        6451 => X"31",  -- 49
        6452 => X"2F",  -- 47
        6453 => X"30",  -- 48
        6454 => X"2E",  -- 46
        6455 => X"2F",  -- 47
        6456 => X"2C",  -- 44
        6457 => X"2C",  -- 44
        6458 => X"2D",  -- 45
        6459 => X"2D",  -- 45
        6460 => X"2B",  -- 43
        6461 => X"2A",  -- 42
        6462 => X"2B",  -- 43
        6463 => X"2E",  -- 46
        6464 => X"30",  -- 48
        6465 => X"30",  -- 48
        6466 => X"31",  -- 49
        6467 => X"34",  -- 52
        6468 => X"39",  -- 57
        6469 => X"40",  -- 64
        6470 => X"48",  -- 72
        6471 => X"4D",  -- 77
        6472 => X"56",  -- 86
        6473 => X"5E",  -- 94
        6474 => X"67",  -- 103
        6475 => X"6C",  -- 108
        6476 => X"6E",  -- 110
        6477 => X"73",  -- 115
        6478 => X"7B",  -- 123
        6479 => X"82",  -- 130
        6480 => X"97",  -- 151
        6481 => X"A5",  -- 165
        6482 => X"A6",  -- 166
        6483 => X"AA",  -- 170
        6484 => X"A4",  -- 164
        6485 => X"9E",  -- 158
        6486 => X"A2",  -- 162
        6487 => X"9A",  -- 154
        6488 => X"93",  -- 147
        6489 => X"9E",  -- 158
        6490 => X"A3",  -- 163
        6491 => X"9F",  -- 159
        6492 => X"9C",  -- 156
        6493 => X"A0",  -- 160
        6494 => X"A3",  -- 163
        6495 => X"9F",  -- 159
        6496 => X"A1",  -- 161
        6497 => X"9B",  -- 155
        6498 => X"A4",  -- 164
        6499 => X"A5",  -- 165
        6500 => X"A3",  -- 163
        6501 => X"9D",  -- 157
        6502 => X"8F",  -- 143
        6503 => X"93",  -- 147
        6504 => X"85",  -- 133
        6505 => X"7D",  -- 125
        6506 => X"7D",  -- 125
        6507 => X"65",  -- 101
        6508 => X"53",  -- 83
        6509 => X"37",  -- 55
        6510 => X"46",  -- 70
        6511 => X"59",  -- 89
        6512 => X"52",  -- 82
        6513 => X"40",  -- 64
        6514 => X"3F",  -- 63
        6515 => X"49",  -- 73
        6516 => X"58",  -- 88
        6517 => X"69",  -- 105
        6518 => X"7C",  -- 124
        6519 => X"83",  -- 131
        6520 => X"82",  -- 130
        6521 => X"87",  -- 135
        6522 => X"8A",  -- 138
        6523 => X"8C",  -- 140
        6524 => X"8B",  -- 139
        6525 => X"8B",  -- 139
        6526 => X"8D",  -- 141
        6527 => X"8F",  -- 143
        6528 => X"88",  -- 136
        6529 => X"8B",  -- 139
        6530 => X"85",  -- 133
        6531 => X"82",  -- 130
        6532 => X"82",  -- 130
        6533 => X"6A",  -- 106
        6534 => X"4F",  -- 79
        6535 => X"4C",  -- 76
        6536 => X"43",  -- 67
        6537 => X"39",  -- 57
        6538 => X"3F",  -- 63
        6539 => X"44",  -- 68
        6540 => X"3C",  -- 60
        6541 => X"43",  -- 67
        6542 => X"50",  -- 80
        6543 => X"4F",  -- 79
        6544 => X"43",  -- 67
        6545 => X"4C",  -- 76
        6546 => X"52",  -- 82
        6547 => X"51",  -- 81
        6548 => X"44",  -- 68
        6549 => X"39",  -- 57
        6550 => X"39",  -- 57
        6551 => X"40",  -- 64
        6552 => X"4C",  -- 76
        6553 => X"50",  -- 80
        6554 => X"55",  -- 85
        6555 => X"58",  -- 88
        6556 => X"5C",  -- 92
        6557 => X"5D",  -- 93
        6558 => X"57",  -- 87
        6559 => X"51",  -- 81
        6560 => X"47",  -- 71
        6561 => X"4D",  -- 77
        6562 => X"5C",  -- 92
        6563 => X"6F",  -- 111
        6564 => X"7A",  -- 122
        6565 => X"74",  -- 116
        6566 => X"63",  -- 99
        6567 => X"54",  -- 84
        6568 => X"3F",  -- 63
        6569 => X"3B",  -- 59
        6570 => X"3B",  -- 59
        6571 => X"46",  -- 70
        6572 => X"55",  -- 85
        6573 => X"5F",  -- 95
        6574 => X"65",  -- 101
        6575 => X"69",  -- 105
        6576 => X"6C",  -- 108
        6577 => X"6A",  -- 106
        6578 => X"68",  -- 104
        6579 => X"69",  -- 105
        6580 => X"6B",  -- 107
        6581 => X"6F",  -- 111
        6582 => X"73",  -- 115
        6583 => X"75",  -- 117
        6584 => X"6D",  -- 109
        6585 => X"6C",  -- 108
        6586 => X"6C",  -- 108
        6587 => X"72",  -- 114
        6588 => X"7B",  -- 123
        6589 => X"82",  -- 130
        6590 => X"83",  -- 131
        6591 => X"83",  -- 131
        6592 => X"81",  -- 129
        6593 => X"7F",  -- 127
        6594 => X"7D",  -- 125
        6595 => X"7D",  -- 125
        6596 => X"82",  -- 130
        6597 => X"87",  -- 135
        6598 => X"8A",  -- 138
        6599 => X"8A",  -- 138
        6600 => X"90",  -- 144
        6601 => X"90",  -- 144
        6602 => X"8F",  -- 143
        6603 => X"8F",  -- 143
        6604 => X"92",  -- 146
        6605 => X"98",  -- 152
        6606 => X"9D",  -- 157
        6607 => X"9F",  -- 159
        6608 => X"A5",  -- 165
        6609 => X"A5",  -- 165
        6610 => X"A6",  -- 166
        6611 => X"A9",  -- 169
        6612 => X"AC",  -- 172
        6613 => X"B1",  -- 177
        6614 => X"B4",  -- 180
        6615 => X"B6",  -- 182
        6616 => X"BA",  -- 186
        6617 => X"BA",  -- 186
        6618 => X"B8",  -- 184
        6619 => X"B6",  -- 182
        6620 => X"B7",  -- 183
        6621 => X"B7",  -- 183
        6622 => X"B0",  -- 176
        6623 => X"A7",  -- 167
        6624 => X"8C",  -- 140
        6625 => X"79",  -- 121
        6626 => X"7C",  -- 124
        6627 => X"8B",  -- 139
        6628 => X"8A",  -- 138
        6629 => X"87",  -- 135
        6630 => X"8B",  -- 139
        6631 => X"91",  -- 145
        6632 => X"90",  -- 144
        6633 => X"95",  -- 149
        6634 => X"96",  -- 150
        6635 => X"97",  -- 151
        6636 => X"98",  -- 152
        6637 => X"9D",  -- 157
        6638 => X"9F",  -- 159
        6639 => X"9E",  -- 158
        6640 => X"A1",  -- 161
        6641 => X"A9",  -- 169
        6642 => X"AF",  -- 175
        6643 => X"B0",  -- 176
        6644 => X"AE",  -- 174
        6645 => X"AD",  -- 173
        6646 => X"AA",  -- 170
        6647 => X"A6",  -- 166
        6648 => X"AD",  -- 173
        6649 => X"AD",  -- 173
        6650 => X"AD",  -- 173
        6651 => X"AE",  -- 174
        6652 => X"AF",  -- 175
        6653 => X"B1",  -- 177
        6654 => X"B3",  -- 179
        6655 => X"B3",  -- 179
        6656 => X"B5",  -- 181
        6657 => X"B3",  -- 179
        6658 => X"B3",  -- 179
        6659 => X"B5",  -- 181
        6660 => X"B6",  -- 182
        6661 => X"B0",  -- 176
        6662 => X"A2",  -- 162
        6663 => X"96",  -- 150
        6664 => X"8D",  -- 141
        6665 => X"7F",  -- 127
        6666 => X"7E",  -- 126
        6667 => X"83",  -- 131
        6668 => X"86",  -- 134
        6669 => X"91",  -- 145
        6670 => X"9C",  -- 156
        6671 => X"98",  -- 152
        6672 => X"97",  -- 151
        6673 => X"9A",  -- 154
        6674 => X"9B",  -- 155
        6675 => X"9C",  -- 156
        6676 => X"9C",  -- 156
        6677 => X"9B",  -- 155
        6678 => X"9C",  -- 156
        6679 => X"9B",  -- 155
        6680 => X"96",  -- 150
        6681 => X"99",  -- 153
        6682 => X"9B",  -- 155
        6683 => X"99",  -- 153
        6684 => X"97",  -- 151
        6685 => X"90",  -- 144
        6686 => X"80",  -- 128
        6687 => X"73",  -- 115
        6688 => X"63",  -- 99
        6689 => X"60",  -- 96
        6690 => X"5F",  -- 95
        6691 => X"5D",  -- 93
        6692 => X"53",  -- 83
        6693 => X"4B",  -- 75
        6694 => X"4A",  -- 74
        6695 => X"51",  -- 81
        6696 => X"72",  -- 114
        6697 => X"8F",  -- 143
        6698 => X"A4",  -- 164
        6699 => X"AD",  -- 173
        6700 => X"B9",  -- 185
        6701 => X"BD",  -- 189
        6702 => X"BC",  -- 188
        6703 => X"C0",  -- 192
        6704 => X"BE",  -- 190
        6705 => X"BE",  -- 190
        6706 => X"BD",  -- 189
        6707 => X"BC",  -- 188
        6708 => X"BC",  -- 188
        6709 => X"BE",  -- 190
        6710 => X"BE",  -- 190
        6711 => X"BE",  -- 190
        6712 => X"C1",  -- 193
        6713 => X"C0",  -- 192
        6714 => X"BD",  -- 189
        6715 => X"B6",  -- 182
        6716 => X"AB",  -- 171
        6717 => X"A3",  -- 163
        6718 => X"A3",  -- 163
        6719 => X"A9",  -- 169
        6720 => X"3D",  -- 61
        6721 => X"3C",  -- 60
        6722 => X"3C",  -- 60
        6723 => X"3B",  -- 59
        6724 => X"3B",  -- 59
        6725 => X"3B",  -- 59
        6726 => X"3B",  -- 59
        6727 => X"3B",  -- 59
        6728 => X"3B",  -- 59
        6729 => X"3C",  -- 60
        6730 => X"3C",  -- 60
        6731 => X"3C",  -- 60
        6732 => X"3D",  -- 61
        6733 => X"3E",  -- 62
        6734 => X"3E",  -- 62
        6735 => X"3E",  -- 62
        6736 => X"3D",  -- 61
        6737 => X"3D",  -- 61
        6738 => X"3D",  -- 61
        6739 => X"3D",  -- 61
        6740 => X"3D",  -- 61
        6741 => X"3D",  -- 61
        6742 => X"3D",  -- 61
        6743 => X"3D",  -- 61
        6744 => X"3D",  -- 61
        6745 => X"3E",  -- 62
        6746 => X"3E",  -- 62
        6747 => X"3F",  -- 63
        6748 => X"3F",  -- 63
        6749 => X"3E",  -- 62
        6750 => X"3E",  -- 62
        6751 => X"3D",  -- 61
        6752 => X"3E",  -- 62
        6753 => X"3C",  -- 60
        6754 => X"3C",  -- 60
        6755 => X"3B",  -- 59
        6756 => X"3A",  -- 58
        6757 => X"39",  -- 57
        6758 => X"38",  -- 56
        6759 => X"37",  -- 55
        6760 => X"34",  -- 52
        6761 => X"34",  -- 52
        6762 => X"34",  -- 52
        6763 => X"33",  -- 51
        6764 => X"33",  -- 51
        6765 => X"33",  -- 51
        6766 => X"33",  -- 51
        6767 => X"33",  -- 51
        6768 => X"32",  -- 50
        6769 => X"32",  -- 50
        6770 => X"31",  -- 49
        6771 => X"30",  -- 48
        6772 => X"30",  -- 48
        6773 => X"2F",  -- 47
        6774 => X"2E",  -- 46
        6775 => X"2E",  -- 46
        6776 => X"2B",  -- 43
        6777 => X"2E",  -- 46
        6778 => X"2E",  -- 46
        6779 => X"2A",  -- 42
        6780 => X"27",  -- 39
        6781 => X"27",  -- 39
        6782 => X"29",  -- 41
        6783 => X"2C",  -- 44
        6784 => X"2F",  -- 47
        6785 => X"31",  -- 49
        6786 => X"33",  -- 51
        6787 => X"39",  -- 57
        6788 => X"3F",  -- 63
        6789 => X"49",  -- 73
        6790 => X"54",  -- 84
        6791 => X"5C",  -- 92
        6792 => X"6A",  -- 106
        6793 => X"73",  -- 115
        6794 => X"7B",  -- 123
        6795 => X"7E",  -- 126
        6796 => X"7D",  -- 125
        6797 => X"7D",  -- 125
        6798 => X"84",  -- 132
        6799 => X"89",  -- 137
        6800 => X"98",  -- 152
        6801 => X"A5",  -- 165
        6802 => X"A9",  -- 169
        6803 => X"AF",  -- 175
        6804 => X"A7",  -- 167
        6805 => X"99",  -- 153
        6806 => X"9A",  -- 154
        6807 => X"95",  -- 149
        6808 => X"97",  -- 151
        6809 => X"9B",  -- 155
        6810 => X"A0",  -- 160
        6811 => X"A1",  -- 161
        6812 => X"A1",  -- 161
        6813 => X"9F",  -- 159
        6814 => X"9F",  -- 159
        6815 => X"9F",  -- 159
        6816 => X"AA",  -- 170
        6817 => X"9F",  -- 159
        6818 => X"A4",  -- 164
        6819 => X"A6",  -- 166
        6820 => X"A4",  -- 164
        6821 => X"9F",  -- 159
        6822 => X"94",  -- 148
        6823 => X"9E",  -- 158
        6824 => X"90",  -- 144
        6825 => X"86",  -- 134
        6826 => X"7E",  -- 126
        6827 => X"62",  -- 98
        6828 => X"54",  -- 84
        6829 => X"42",  -- 66
        6830 => X"4F",  -- 79
        6831 => X"5B",  -- 91
        6832 => X"4E",  -- 78
        6833 => X"40",  -- 64
        6834 => X"49",  -- 73
        6835 => X"55",  -- 85
        6836 => X"63",  -- 99
        6837 => X"65",  -- 101
        6838 => X"7B",  -- 123
        6839 => X"84",  -- 132
        6840 => X"81",  -- 129
        6841 => X"85",  -- 133
        6842 => X"87",  -- 135
        6843 => X"88",  -- 136
        6844 => X"86",  -- 134
        6845 => X"85",  -- 133
        6846 => X"86",  -- 134
        6847 => X"87",  -- 135
        6848 => X"85",  -- 133
        6849 => X"84",  -- 132
        6850 => X"7F",  -- 127
        6851 => X"7B",  -- 123
        6852 => X"77",  -- 119
        6853 => X"67",  -- 103
        6854 => X"52",  -- 82
        6855 => X"4A",  -- 74
        6856 => X"37",  -- 55
        6857 => X"42",  -- 66
        6858 => X"52",  -- 82
        6859 => X"57",  -- 87
        6860 => X"4E",  -- 78
        6861 => X"46",  -- 70
        6862 => X"40",  -- 64
        6863 => X"37",  -- 55
        6864 => X"41",  -- 65
        6865 => X"49",  -- 73
        6866 => X"49",  -- 73
        6867 => X"3A",  -- 58
        6868 => X"2F",  -- 47
        6869 => X"2F",  -- 47
        6870 => X"37",  -- 55
        6871 => X"39",  -- 57
        6872 => X"42",  -- 66
        6873 => X"47",  -- 71
        6874 => X"4F",  -- 79
        6875 => X"54",  -- 84
        6876 => X"58",  -- 88
        6877 => X"53",  -- 83
        6878 => X"46",  -- 70
        6879 => X"39",  -- 57
        6880 => X"31",  -- 49
        6881 => X"34",  -- 52
        6882 => X"43",  -- 67
        6883 => X"59",  -- 89
        6884 => X"68",  -- 104
        6885 => X"64",  -- 100
        6886 => X"53",  -- 83
        6887 => X"46",  -- 70
        6888 => X"42",  -- 66
        6889 => X"42",  -- 66
        6890 => X"47",  -- 71
        6891 => X"4E",  -- 78
        6892 => X"54",  -- 84
        6893 => X"58",  -- 88
        6894 => X"5E",  -- 94
        6895 => X"65",  -- 101
        6896 => X"6A",  -- 106
        6897 => X"6A",  -- 106
        6898 => X"6B",  -- 107
        6899 => X"6E",  -- 110
        6900 => X"72",  -- 114
        6901 => X"73",  -- 115
        6902 => X"73",  -- 115
        6903 => X"74",  -- 116
        6904 => X"6E",  -- 110
        6905 => X"6D",  -- 109
        6906 => X"6E",  -- 110
        6907 => X"75",  -- 117
        6908 => X"7E",  -- 126
        6909 => X"82",  -- 130
        6910 => X"7F",  -- 127
        6911 => X"7B",  -- 123
        6912 => X"7A",  -- 122
        6913 => X"7A",  -- 122
        6914 => X"79",  -- 121
        6915 => X"79",  -- 121
        6916 => X"7F",  -- 127
        6917 => X"88",  -- 136
        6918 => X"8D",  -- 141
        6919 => X"8E",  -- 142
        6920 => X"8A",  -- 138
        6921 => X"8A",  -- 138
        6922 => X"8A",  -- 138
        6923 => X"8A",  -- 138
        6924 => X"91",  -- 145
        6925 => X"99",  -- 153
        6926 => X"9F",  -- 159
        6927 => X"A0",  -- 160
        6928 => X"A2",  -- 162
        6929 => X"A3",  -- 163
        6930 => X"A4",  -- 164
        6931 => X"A7",  -- 167
        6932 => X"AA",  -- 170
        6933 => X"AE",  -- 174
        6934 => X"B3",  -- 179
        6935 => X"B4",  -- 180
        6936 => X"B5",  -- 181
        6937 => X"B7",  -- 183
        6938 => X"B6",  -- 182
        6939 => X"B5",  -- 181
        6940 => X"B7",  -- 183
        6941 => X"B8",  -- 184
        6942 => X"B2",  -- 178
        6943 => X"AA",  -- 170
        6944 => X"97",  -- 151
        6945 => X"85",  -- 133
        6946 => X"83",  -- 131
        6947 => X"8B",  -- 139
        6948 => X"86",  -- 134
        6949 => X"81",  -- 129
        6950 => X"87",  -- 135
        6951 => X"8C",  -- 140
        6952 => X"91",  -- 145
        6953 => X"93",  -- 147
        6954 => X"93",  -- 147
        6955 => X"94",  -- 148
        6956 => X"95",  -- 149
        6957 => X"9A",  -- 154
        6958 => X"9D",  -- 157
        6959 => X"9B",  -- 155
        6960 => X"A5",  -- 165
        6961 => X"AD",  -- 173
        6962 => X"B2",  -- 178
        6963 => X"B1",  -- 177
        6964 => X"AE",  -- 174
        6965 => X"AB",  -- 171
        6966 => X"A8",  -- 168
        6967 => X"A5",  -- 165
        6968 => X"AC",  -- 172
        6969 => X"AB",  -- 171
        6970 => X"AA",  -- 170
        6971 => X"AA",  -- 170
        6972 => X"AC",  -- 172
        6973 => X"AE",  -- 174
        6974 => X"B2",  -- 178
        6975 => X"B3",  -- 179
        6976 => X"B4",  -- 180
        6977 => X"B3",  -- 179
        6978 => X"B4",  -- 180
        6979 => X"B5",  -- 181
        6980 => X"B5",  -- 181
        6981 => X"B0",  -- 176
        6982 => X"A5",  -- 165
        6983 => X"9B",  -- 155
        6984 => X"8D",  -- 141
        6985 => X"80",  -- 128
        6986 => X"73",  -- 115
        6987 => X"73",  -- 115
        6988 => X"7E",  -- 126
        6989 => X"8A",  -- 138
        6990 => X"91",  -- 145
        6991 => X"97",  -- 151
        6992 => X"99",  -- 153
        6993 => X"9E",  -- 158
        6994 => X"A0",  -- 160
        6995 => X"A2",  -- 162
        6996 => X"A2",  -- 162
        6997 => X"9E",  -- 158
        6998 => X"9C",  -- 156
        6999 => X"9B",  -- 155
        7000 => X"99",  -- 153
        7001 => X"9A",  -- 154
        7002 => X"9A",  -- 154
        7003 => X"9C",  -- 156
        7004 => X"9E",  -- 158
        7005 => X"9D",  -- 157
        7006 => X"96",  -- 150
        7007 => X"8E",  -- 142
        7008 => X"78",  -- 120
        7009 => X"69",  -- 105
        7010 => X"5C",  -- 92
        7011 => X"5B",  -- 91
        7012 => X"59",  -- 89
        7013 => X"54",  -- 84
        7014 => X"55",  -- 85
        7015 => X"5C",  -- 92
        7016 => X"71",  -- 113
        7017 => X"8C",  -- 140
        7018 => X"A1",  -- 161
        7019 => X"AA",  -- 170
        7020 => X"B7",  -- 183
        7021 => X"BB",  -- 187
        7022 => X"BB",  -- 187
        7023 => X"BB",  -- 187
        7024 => X"C0",  -- 192
        7025 => X"C0",  -- 192
        7026 => X"C0",  -- 192
        7027 => X"C2",  -- 194
        7028 => X"C3",  -- 195
        7029 => X"C2",  -- 194
        7030 => X"C4",  -- 196
        7031 => X"C3",  -- 195
        7032 => X"BF",  -- 191
        7033 => X"C0",  -- 192
        7034 => X"BF",  -- 191
        7035 => X"B9",  -- 185
        7036 => X"AC",  -- 172
        7037 => X"A3",  -- 163
        7038 => X"A3",  -- 163
        7039 => X"A6",  -- 166
        7040 => X"3D",  -- 61
        7041 => X"3C",  -- 60
        7042 => X"3B",  -- 59
        7043 => X"3B",  -- 59
        7044 => X"3B",  -- 59
        7045 => X"3B",  -- 59
        7046 => X"3B",  -- 59
        7047 => X"3C",  -- 60
        7048 => X"3C",  -- 60
        7049 => X"3C",  -- 60
        7050 => X"3C",  -- 60
        7051 => X"3D",  -- 61
        7052 => X"3D",  -- 61
        7053 => X"3E",  -- 62
        7054 => X"3E",  -- 62
        7055 => X"3E",  -- 62
        7056 => X"3D",  -- 61
        7057 => X"3D",  -- 61
        7058 => X"3D",  -- 61
        7059 => X"3D",  -- 61
        7060 => X"3D",  -- 61
        7061 => X"3D",  -- 61
        7062 => X"3D",  -- 61
        7063 => X"3D",  -- 61
        7064 => X"3D",  -- 61
        7065 => X"3E",  -- 62
        7066 => X"3E",  -- 62
        7067 => X"3E",  -- 62
        7068 => X"3E",  -- 62
        7069 => X"3E",  -- 62
        7070 => X"3D",  -- 61
        7071 => X"3D",  -- 61
        7072 => X"3E",  -- 62
        7073 => X"3C",  -- 60
        7074 => X"3C",  -- 60
        7075 => X"3B",  -- 59
        7076 => X"3A",  -- 58
        7077 => X"38",  -- 56
        7078 => X"37",  -- 55
        7079 => X"37",  -- 55
        7080 => X"34",  -- 52
        7081 => X"34",  -- 52
        7082 => X"34",  -- 52
        7083 => X"34",  -- 52
        7084 => X"34",  -- 52
        7085 => X"34",  -- 52
        7086 => X"34",  -- 52
        7087 => X"34",  -- 52
        7088 => X"32",  -- 50
        7089 => X"32",  -- 50
        7090 => X"31",  -- 49
        7091 => X"31",  -- 49
        7092 => X"30",  -- 48
        7093 => X"30",  -- 48
        7094 => X"2F",  -- 47
        7095 => X"2E",  -- 46
        7096 => X"2B",  -- 43
        7097 => X"2C",  -- 44
        7098 => X"2C",  -- 44
        7099 => X"2A",  -- 42
        7100 => X"29",  -- 41
        7101 => X"2B",  -- 43
        7102 => X"31",  -- 49
        7103 => X"36",  -- 54
        7104 => X"3C",  -- 60
        7105 => X"3E",  -- 62
        7106 => X"44",  -- 68
        7107 => X"4A",  -- 74
        7108 => X"52",  -- 82
        7109 => X"5C",  -- 92
        7110 => X"65",  -- 101
        7111 => X"6B",  -- 107
        7112 => X"78",  -- 120
        7113 => X"81",  -- 129
        7114 => X"88",  -- 136
        7115 => X"87",  -- 135
        7116 => X"83",  -- 131
        7117 => X"84",  -- 132
        7118 => X"8A",  -- 138
        7119 => X"91",  -- 145
        7120 => X"9F",  -- 159
        7121 => X"A4",  -- 164
        7122 => X"A2",  -- 162
        7123 => X"AD",  -- 173
        7124 => X"A7",  -- 167
        7125 => X"95",  -- 149
        7126 => X"96",  -- 150
        7127 => X"93",  -- 147
        7128 => X"9C",  -- 156
        7129 => X"98",  -- 152
        7130 => X"9B",  -- 155
        7131 => X"A3",  -- 163
        7132 => X"A4",  -- 164
        7133 => X"9C",  -- 156
        7134 => X"99",  -- 153
        7135 => X"9D",  -- 157
        7136 => X"A7",  -- 167
        7137 => X"9F",  -- 159
        7138 => X"A5",  -- 165
        7139 => X"A0",  -- 160
        7140 => X"9D",  -- 157
        7141 => X"A0",  -- 160
        7142 => X"99",  -- 153
        7143 => X"9E",  -- 158
        7144 => X"93",  -- 147
        7145 => X"86",  -- 134
        7146 => X"7A",  -- 122
        7147 => X"60",  -- 96
        7148 => X"60",  -- 96
        7149 => X"5A",  -- 90
        7150 => X"61",  -- 97
        7151 => X"5C",  -- 92
        7152 => X"57",  -- 87
        7153 => X"55",  -- 85
        7154 => X"6A",  -- 106
        7155 => X"6D",  -- 109
        7156 => X"74",  -- 116
        7157 => X"6F",  -- 111
        7158 => X"83",  -- 131
        7159 => X"89",  -- 137
        7160 => X"80",  -- 128
        7161 => X"82",  -- 130
        7162 => X"87",  -- 135
        7163 => X"87",  -- 135
        7164 => X"87",  -- 135
        7165 => X"85",  -- 133
        7166 => X"82",  -- 130
        7167 => X"81",  -- 129
        7168 => X"82",  -- 130
        7169 => X"7E",  -- 126
        7170 => X"7D",  -- 125
        7171 => X"79",  -- 121
        7172 => X"6F",  -- 111
        7173 => X"69",  -- 105
        7174 => X"5F",  -- 95
        7175 => X"50",  -- 80
        7176 => X"41",  -- 65
        7177 => X"54",  -- 84
        7178 => X"66",  -- 102
        7179 => X"6B",  -- 107
        7180 => X"62",  -- 98
        7181 => X"4E",  -- 78
        7182 => X"3D",  -- 61
        7183 => X"3B",  -- 59
        7184 => X"51",  -- 81
        7185 => X"4F",  -- 79
        7186 => X"44",  -- 68
        7187 => X"38",  -- 56
        7188 => X"32",  -- 50
        7189 => X"32",  -- 50
        7190 => X"33",  -- 51
        7191 => X"2F",  -- 47
        7192 => X"2D",  -- 45
        7193 => X"33",  -- 51
        7194 => X"3B",  -- 59
        7195 => X"3F",  -- 63
        7196 => X"3D",  -- 61
        7197 => X"38",  -- 56
        7198 => X"2D",  -- 45
        7199 => X"23",  -- 35
        7200 => X"31",  -- 49
        7201 => X"30",  -- 48
        7202 => X"3B",  -- 59
        7203 => X"4F",  -- 79
        7204 => X"5E",  -- 94
        7205 => X"5A",  -- 90
        7206 => X"4C",  -- 76
        7207 => X"40",  -- 64
        7208 => X"3D",  -- 61
        7209 => X"40",  -- 64
        7210 => X"48",  -- 72
        7211 => X"4F",  -- 79
        7212 => X"50",  -- 80
        7213 => X"51",  -- 81
        7214 => X"57",  -- 87
        7215 => X"5F",  -- 95
        7216 => X"6B",  -- 107
        7217 => X"6B",  -- 107
        7218 => X"6E",  -- 110
        7219 => X"73",  -- 115
        7220 => X"78",  -- 120
        7221 => X"77",  -- 119
        7222 => X"73",  -- 115
        7223 => X"70",  -- 112
        7224 => X"73",  -- 115
        7225 => X"74",  -- 116
        7226 => X"76",  -- 118
        7227 => X"79",  -- 121
        7228 => X"79",  -- 121
        7229 => X"77",  -- 119
        7230 => X"73",  -- 115
        7231 => X"6F",  -- 111
        7232 => X"7E",  -- 126
        7233 => X"7F",  -- 127
        7234 => X"7D",  -- 125
        7235 => X"78",  -- 120
        7236 => X"79",  -- 121
        7237 => X"7F",  -- 127
        7238 => X"84",  -- 132
        7239 => X"84",  -- 132
        7240 => X"85",  -- 133
        7241 => X"8B",  -- 139
        7242 => X"8D",  -- 141
        7243 => X"8D",  -- 141
        7244 => X"8F",  -- 143
        7245 => X"96",  -- 150
        7246 => X"9B",  -- 155
        7247 => X"9D",  -- 157
        7248 => X"9D",  -- 157
        7249 => X"9E",  -- 158
        7250 => X"A0",  -- 160
        7251 => X"A4",  -- 164
        7252 => X"A8",  -- 168
        7253 => X"AC",  -- 172
        7254 => X"B0",  -- 176
        7255 => X"B3",  -- 179
        7256 => X"B1",  -- 177
        7257 => X"B4",  -- 180
        7258 => X"B7",  -- 183
        7259 => X"B8",  -- 184
        7260 => X"B8",  -- 184
        7261 => X"B9",  -- 185
        7262 => X"B4",  -- 180
        7263 => X"AF",  -- 175
        7264 => X"A5",  -- 165
        7265 => X"94",  -- 148
        7266 => X"8D",  -- 141
        7267 => X"8C",  -- 140
        7268 => X"85",  -- 133
        7269 => X"82",  -- 130
        7270 => X"88",  -- 136
        7271 => X"8A",  -- 138
        7272 => X"90",  -- 144
        7273 => X"92",  -- 146
        7274 => X"90",  -- 144
        7275 => X"91",  -- 145
        7276 => X"93",  -- 147
        7277 => X"9A",  -- 154
        7278 => X"9D",  -- 157
        7279 => X"9D",  -- 157
        7280 => X"A5",  -- 165
        7281 => X"AC",  -- 172
        7282 => X"B1",  -- 177
        7283 => X"AE",  -- 174
        7284 => X"AA",  -- 170
        7285 => X"A8",  -- 168
        7286 => X"A7",  -- 167
        7287 => X"A4",  -- 164
        7288 => X"A7",  -- 167
        7289 => X"A7",  -- 167
        7290 => X"A9",  -- 169
        7291 => X"AB",  -- 171
        7292 => X"AD",  -- 173
        7293 => X"B0",  -- 176
        7294 => X"B3",  -- 179
        7295 => X"B6",  -- 182
        7296 => X"B1",  -- 177
        7297 => X"B2",  -- 178
        7298 => X"B4",  -- 180
        7299 => X"B7",  -- 183
        7300 => X"B5",  -- 181
        7301 => X"B2",  -- 178
        7302 => X"AB",  -- 171
        7303 => X"A5",  -- 165
        7304 => X"93",  -- 147
        7305 => X"8D",  -- 141
        7306 => X"72",  -- 114
        7307 => X"68",  -- 104
        7308 => X"76",  -- 118
        7309 => X"78",  -- 120
        7310 => X"78",  -- 120
        7311 => X"8A",  -- 138
        7312 => X"9C",  -- 156
        7313 => X"9F",  -- 159
        7314 => X"A2",  -- 162
        7315 => X"A4",  -- 164
        7316 => X"A3",  -- 163
        7317 => X"9E",  -- 158
        7318 => X"9B",  -- 155
        7319 => X"99",  -- 153
        7320 => X"99",  -- 153
        7321 => X"9B",  -- 155
        7322 => X"9B",  -- 155
        7323 => X"9C",  -- 156
        7324 => X"A1",  -- 161
        7325 => X"A2",  -- 162
        7326 => X"9D",  -- 157
        7327 => X"96",  -- 150
        7328 => X"83",  -- 131
        7329 => X"6F",  -- 111
        7330 => X"61",  -- 97
        7331 => X"63",  -- 99
        7332 => X"64",  -- 100
        7333 => X"5D",  -- 93
        7334 => X"5A",  -- 90
        7335 => X"5C",  -- 92
        7336 => X"69",  -- 105
        7337 => X"84",  -- 132
        7338 => X"97",  -- 151
        7339 => X"A4",  -- 164
        7340 => X"B0",  -- 176
        7341 => X"B5",  -- 181
        7342 => X"B5",  -- 181
        7343 => X"B7",  -- 183
        7344 => X"BE",  -- 190
        7345 => X"BE",  -- 190
        7346 => X"BE",  -- 190
        7347 => X"BE",  -- 190
        7348 => X"C0",  -- 192
        7349 => X"C0",  -- 192
        7350 => X"C2",  -- 194
        7351 => X"C2",  -- 194
        7352 => X"BC",  -- 188
        7353 => X"BF",  -- 191
        7354 => X"BF",  -- 191
        7355 => X"B8",  -- 184
        7356 => X"AC",  -- 172
        7357 => X"A5",  -- 165
        7358 => X"A6",  -- 166
        7359 => X"AA",  -- 170
        7360 => X"3C",  -- 60
        7361 => X"3C",  -- 60
        7362 => X"3B",  -- 59
        7363 => X"3B",  -- 59
        7364 => X"3B",  -- 59
        7365 => X"3B",  -- 59
        7366 => X"3C",  -- 60
        7367 => X"3C",  -- 60
        7368 => X"3C",  -- 60
        7369 => X"3C",  -- 60
        7370 => X"3C",  -- 60
        7371 => X"3D",  -- 61
        7372 => X"3D",  -- 61
        7373 => X"3E",  -- 62
        7374 => X"3E",  -- 62
        7375 => X"3F",  -- 63
        7376 => X"3D",  -- 61
        7377 => X"3D",  -- 61
        7378 => X"3D",  -- 61
        7379 => X"3D",  -- 61
        7380 => X"3D",  -- 61
        7381 => X"3D",  -- 61
        7382 => X"3D",  -- 61
        7383 => X"3D",  -- 61
        7384 => X"3D",  -- 61
        7385 => X"3E",  -- 62
        7386 => X"3E",  -- 62
        7387 => X"3E",  -- 62
        7388 => X"3E",  -- 62
        7389 => X"3E",  -- 62
        7390 => X"3D",  -- 61
        7391 => X"3C",  -- 60
        7392 => X"3E",  -- 62
        7393 => X"3C",  -- 60
        7394 => X"3C",  -- 60
        7395 => X"3B",  -- 59
        7396 => X"39",  -- 57
        7397 => X"38",  -- 56
        7398 => X"37",  -- 55
        7399 => X"37",  -- 55
        7400 => X"33",  -- 51
        7401 => X"33",  -- 51
        7402 => X"34",  -- 52
        7403 => X"34",  -- 52
        7404 => X"34",  -- 52
        7405 => X"34",  -- 52
        7406 => X"34",  -- 52
        7407 => X"34",  -- 52
        7408 => X"32",  -- 50
        7409 => X"32",  -- 50
        7410 => X"32",  -- 50
        7411 => X"32",  -- 50
        7412 => X"31",  -- 49
        7413 => X"30",  -- 48
        7414 => X"30",  -- 48
        7415 => X"2F",  -- 47
        7416 => X"2E",  -- 46
        7417 => X"2F",  -- 47
        7418 => X"31",  -- 49
        7419 => X"32",  -- 50
        7420 => X"32",  -- 50
        7421 => X"36",  -- 54
        7422 => X"3F",  -- 63
        7423 => X"45",  -- 69
        7424 => X"50",  -- 80
        7425 => X"54",  -- 84
        7426 => X"5C",  -- 92
        7427 => X"62",  -- 98
        7428 => X"6A",  -- 106
        7429 => X"70",  -- 112
        7430 => X"76",  -- 118
        7431 => X"79",  -- 121
        7432 => X"7E",  -- 126
        7433 => X"84",  -- 132
        7434 => X"8A",  -- 138
        7435 => X"89",  -- 137
        7436 => X"86",  -- 134
        7437 => X"88",  -- 136
        7438 => X"91",  -- 145
        7439 => X"9A",  -- 154
        7440 => X"A8",  -- 168
        7441 => X"A4",  -- 164
        7442 => X"9C",  -- 156
        7443 => X"A6",  -- 166
        7444 => X"A2",  -- 162
        7445 => X"93",  -- 147
        7446 => X"96",  -- 150
        7447 => X"98",  -- 152
        7448 => X"A2",  -- 162
        7449 => X"97",  -- 151
        7450 => X"99",  -- 153
        7451 => X"A4",  -- 164
        7452 => X"A4",  -- 164
        7453 => X"99",  -- 153
        7454 => X"95",  -- 149
        7455 => X"9B",  -- 155
        7456 => X"9C",  -- 156
        7457 => X"9E",  -- 158
        7458 => X"A4",  -- 164
        7459 => X"9A",  -- 154
        7460 => X"99",  -- 153
        7461 => X"A1",  -- 161
        7462 => X"98",  -- 152
        7463 => X"96",  -- 150
        7464 => X"8F",  -- 143
        7465 => X"82",  -- 130
        7466 => X"76",  -- 118
        7467 => X"63",  -- 99
        7468 => X"71",  -- 113
        7469 => X"71",  -- 113
        7470 => X"70",  -- 112
        7471 => X"5D",  -- 93
        7472 => X"71",  -- 113
        7473 => X"79",  -- 121
        7474 => X"8F",  -- 143
        7475 => X"85",  -- 133
        7476 => X"83",  -- 131
        7477 => X"7B",  -- 123
        7478 => X"8D",  -- 141
        7479 => X"8B",  -- 139
        7480 => X"7C",  -- 124
        7481 => X"80",  -- 128
        7482 => X"86",  -- 134
        7483 => X"89",  -- 137
        7484 => X"8C",  -- 140
        7485 => X"89",  -- 137
        7486 => X"85",  -- 133
        7487 => X"82",  -- 130
        7488 => X"7F",  -- 127
        7489 => X"7A",  -- 122
        7490 => X"80",  -- 128
        7491 => X"7D",  -- 125
        7492 => X"6F",  -- 111
        7493 => X"6E",  -- 110
        7494 => X"6B",  -- 107
        7495 => X"56",  -- 86
        7496 => X"61",  -- 97
        7497 => X"6D",  -- 109
        7498 => X"6E",  -- 110
        7499 => X"6C",  -- 108
        7500 => X"67",  -- 103
        7501 => X"53",  -- 83
        7502 => X"4F",  -- 79
        7503 => X"63",  -- 99
        7504 => X"67",  -- 103
        7505 => X"5B",  -- 91
        7506 => X"4E",  -- 78
        7507 => X"48",  -- 72
        7508 => X"44",  -- 68
        7509 => X"3E",  -- 62
        7510 => X"33",  -- 51
        7511 => X"29",  -- 41
        7512 => X"35",  -- 53
        7513 => X"35",  -- 53
        7514 => X"30",  -- 48
        7515 => X"28",  -- 40
        7516 => X"25",  -- 37
        7517 => X"2A",  -- 42
        7518 => X"32",  -- 50
        7519 => X"36",  -- 54
        7520 => X"34",  -- 52
        7521 => X"31",  -- 49
        7522 => X"36",  -- 54
        7523 => X"45",  -- 69
        7524 => X"50",  -- 80
        7525 => X"4C",  -- 76
        7526 => X"40",  -- 64
        7527 => X"35",  -- 53
        7528 => X"32",  -- 50
        7529 => X"38",  -- 56
        7530 => X"41",  -- 65
        7531 => X"4B",  -- 75
        7532 => X"4E",  -- 78
        7533 => X"4F",  -- 79
        7534 => X"55",  -- 85
        7535 => X"5D",  -- 93
        7536 => X"68",  -- 104
        7537 => X"6A",  -- 106
        7538 => X"6C",  -- 108
        7539 => X"70",  -- 112
        7540 => X"73",  -- 115
        7541 => X"74",  -- 116
        7542 => X"70",  -- 112
        7543 => X"6C",  -- 108
        7544 => X"70",  -- 112
        7545 => X"74",  -- 116
        7546 => X"78",  -- 120
        7547 => X"79",  -- 121
        7548 => X"76",  -- 118
        7549 => X"72",  -- 114
        7550 => X"70",  -- 112
        7551 => X"6F",  -- 111
        7552 => X"7E",  -- 126
        7553 => X"80",  -- 128
        7554 => X"7E",  -- 126
        7555 => X"76",  -- 118
        7556 => X"74",  -- 116
        7557 => X"78",  -- 120
        7558 => X"7C",  -- 124
        7559 => X"7C",  -- 124
        7560 => X"84",  -- 132
        7561 => X"8E",  -- 142
        7562 => X"94",  -- 148
        7563 => X"92",  -- 146
        7564 => X"8F",  -- 143
        7565 => X"92",  -- 146
        7566 => X"95",  -- 149
        7567 => X"97",  -- 151
        7568 => X"98",  -- 152
        7569 => X"99",  -- 153
        7570 => X"9D",  -- 157
        7571 => X"A2",  -- 162
        7572 => X"A7",  -- 167
        7573 => X"AB",  -- 171
        7574 => X"AF",  -- 175
        7575 => X"B1",  -- 177
        7576 => X"B2",  -- 178
        7577 => X"B5",  -- 181
        7578 => X"B9",  -- 185
        7579 => X"BA",  -- 186
        7580 => X"BB",  -- 187
        7581 => X"BC",  -- 188
        7582 => X"B8",  -- 184
        7583 => X"B3",  -- 179
        7584 => X"AA",  -- 170
        7585 => X"9A",  -- 154
        7586 => X"90",  -- 144
        7587 => X"8B",  -- 139
        7588 => X"82",  -- 130
        7589 => X"81",  -- 129
        7590 => X"88",  -- 136
        7591 => X"89",  -- 137
        7592 => X"90",  -- 144
        7593 => X"91",  -- 145
        7594 => X"8F",  -- 143
        7595 => X"8E",  -- 142
        7596 => X"93",  -- 147
        7597 => X"9B",  -- 155
        7598 => X"9F",  -- 159
        7599 => X"9F",  -- 159
        7600 => X"A4",  -- 164
        7601 => X"AB",  -- 171
        7602 => X"B0",  -- 176
        7603 => X"AE",  -- 174
        7604 => X"AB",  -- 171
        7605 => X"AA",  -- 170
        7606 => X"AB",  -- 171
        7607 => X"AA",  -- 170
        7608 => X"A3",  -- 163
        7609 => X"A5",  -- 165
        7610 => X"A9",  -- 169
        7611 => X"AC",  -- 172
        7612 => X"AF",  -- 175
        7613 => X"B3",  -- 179
        7614 => X"B5",  -- 181
        7615 => X"B8",  -- 184
        7616 => X"AF",  -- 175
        7617 => X"B2",  -- 178
        7618 => X"B5",  -- 181
        7619 => X"B8",  -- 184
        7620 => X"B6",  -- 182
        7621 => X"B5",  -- 181
        7622 => X"B1",  -- 177
        7623 => X"AE",  -- 174
        7624 => X"9B",  -- 155
        7625 => X"9A",  -- 154
        7626 => X"79",  -- 121
        7627 => X"66",  -- 102
        7628 => X"71",  -- 113
        7629 => X"6A",  -- 106
        7630 => X"63",  -- 99
        7631 => X"7C",  -- 124
        7632 => X"94",  -- 148
        7633 => X"97",  -- 151
        7634 => X"9E",  -- 158
        7635 => X"A0",  -- 160
        7636 => X"A2",  -- 162
        7637 => X"A2",  -- 162
        7638 => X"A0",  -- 160
        7639 => X"A1",  -- 161
        7640 => X"99",  -- 153
        7641 => X"9D",  -- 157
        7642 => X"A0",  -- 160
        7643 => X"A3",  -- 163
        7644 => X"A5",  -- 165
        7645 => X"A5",  -- 165
        7646 => X"9A",  -- 154
        7647 => X"91",  -- 145
        7648 => X"8B",  -- 139
        7649 => X"7C",  -- 124
        7650 => X"75",  -- 117
        7651 => X"76",  -- 118
        7652 => X"6B",  -- 107
        7653 => X"56",  -- 86
        7654 => X"4B",  -- 75
        7655 => X"4E",  -- 78
        7656 => X"55",  -- 85
        7657 => X"70",  -- 112
        7658 => X"88",  -- 136
        7659 => X"99",  -- 153
        7660 => X"AB",  -- 171
        7661 => X"B5",  -- 181
        7662 => X"B7",  -- 183
        7663 => X"BB",  -- 187
        7664 => X"BD",  -- 189
        7665 => X"BB",  -- 187
        7666 => X"B9",  -- 185
        7667 => X"B7",  -- 183
        7668 => X"B7",  -- 183
        7669 => X"B9",  -- 185
        7670 => X"BB",  -- 187
        7671 => X"BC",  -- 188
        7672 => X"BB",  -- 187
        7673 => X"BE",  -- 190
        7674 => X"BF",  -- 191
        7675 => X"B7",  -- 183
        7676 => X"AB",  -- 171
        7677 => X"A6",  -- 166
        7678 => X"A8",  -- 168
        7679 => X"AD",  -- 173
        7680 => X"3D",  -- 61
        7681 => X"3D",  -- 61
        7682 => X"3C",  -- 60
        7683 => X"3C",  -- 60
        7684 => X"3D",  -- 61
        7685 => X"3D",  -- 61
        7686 => X"3E",  -- 62
        7687 => X"3F",  -- 63
        7688 => X"3E",  -- 62
        7689 => X"3E",  -- 62
        7690 => X"3F",  -- 63
        7691 => X"3F",  -- 63
        7692 => X"3F",  -- 63
        7693 => X"3F",  -- 63
        7694 => X"3E",  -- 62
        7695 => X"3E",  -- 62
        7696 => X"3E",  -- 62
        7697 => X"3E",  -- 62
        7698 => X"3E",  -- 62
        7699 => X"3E",  -- 62
        7700 => X"3D",  -- 61
        7701 => X"3D",  -- 61
        7702 => X"3D",  -- 61
        7703 => X"3D",  -- 61
        7704 => X"3F",  -- 63
        7705 => X"3E",  -- 62
        7706 => X"3E",  -- 62
        7707 => X"3E",  -- 62
        7708 => X"3E",  -- 62
        7709 => X"3D",  -- 61
        7710 => X"3D",  -- 61
        7711 => X"3D",  -- 61
        7712 => X"3C",  -- 60
        7713 => X"3C",  -- 60
        7714 => X"3C",  -- 60
        7715 => X"3C",  -- 60
        7716 => X"3B",  -- 59
        7717 => X"39",  -- 57
        7718 => X"38",  -- 56
        7719 => X"36",  -- 54
        7720 => X"36",  -- 54
        7721 => X"34",  -- 52
        7722 => X"31",  -- 49
        7723 => X"31",  -- 49
        7724 => X"32",  -- 50
        7725 => X"33",  -- 51
        7726 => X"33",  -- 51
        7727 => X"33",  -- 51
        7728 => X"33",  -- 51
        7729 => X"34",  -- 52
        7730 => X"33",  -- 51
        7731 => X"30",  -- 48
        7732 => X"2F",  -- 47
        7733 => X"2E",  -- 46
        7734 => X"2E",  -- 46
        7735 => X"2F",  -- 47
        7736 => X"35",  -- 53
        7737 => X"3C",  -- 60
        7738 => X"43",  -- 67
        7739 => X"49",  -- 73
        7740 => X"4A",  -- 74
        7741 => X"50",  -- 80
        7742 => X"5B",  -- 91
        7743 => X"62",  -- 98
        7744 => X"6B",  -- 107
        7745 => X"6D",  -- 109
        7746 => X"72",  -- 114
        7747 => X"76",  -- 118
        7748 => X"7D",  -- 125
        7749 => X"7F",  -- 127
        7750 => X"7E",  -- 126
        7751 => X"7E",  -- 126
        7752 => X"7F",  -- 127
        7753 => X"85",  -- 133
        7754 => X"81",  -- 129
        7755 => X"80",  -- 128
        7756 => X"8B",  -- 139
        7757 => X"96",  -- 150
        7758 => X"9E",  -- 158
        7759 => X"A9",  -- 169
        7760 => X"A8",  -- 168
        7761 => X"A2",  -- 162
        7762 => X"A2",  -- 162
        7763 => X"95",  -- 149
        7764 => X"9E",  -- 158
        7765 => X"9D",  -- 157
        7766 => X"A1",  -- 161
        7767 => X"97",  -- 151
        7768 => X"A0",  -- 160
        7769 => X"8E",  -- 142
        7770 => X"95",  -- 149
        7771 => X"99",  -- 153
        7772 => X"A9",  -- 169
        7773 => X"96",  -- 150
        7774 => X"92",  -- 146
        7775 => X"8D",  -- 141
        7776 => X"98",  -- 152
        7777 => X"9E",  -- 158
        7778 => X"9E",  -- 158
        7779 => X"A1",  -- 161
        7780 => X"99",  -- 153
        7781 => X"98",  -- 152
        7782 => X"A2",  -- 162
        7783 => X"97",  -- 151
        7784 => X"93",  -- 147
        7785 => X"77",  -- 119
        7786 => X"6C",  -- 108
        7787 => X"7B",  -- 123
        7788 => X"7A",  -- 122
        7789 => X"8D",  -- 141
        7790 => X"7C",  -- 124
        7791 => X"7C",  -- 124
        7792 => X"8E",  -- 142
        7793 => X"91",  -- 145
        7794 => X"95",  -- 149
        7795 => X"99",  -- 153
        7796 => X"8B",  -- 139
        7797 => X"76",  -- 118
        7798 => X"9C",  -- 156
        7799 => X"84",  -- 132
        7800 => X"80",  -- 128
        7801 => X"8C",  -- 140
        7802 => X"85",  -- 133
        7803 => X"8A",  -- 138
        7804 => X"8F",  -- 143
        7805 => X"86",  -- 134
        7806 => X"83",  -- 131
        7807 => X"7C",  -- 124
        7808 => X"73",  -- 115
        7809 => X"73",  -- 115
        7810 => X"72",  -- 114
        7811 => X"77",  -- 119
        7812 => X"79",  -- 121
        7813 => X"6E",  -- 110
        7814 => X"6A",  -- 106
        7815 => X"74",  -- 116
        7816 => X"77",  -- 119
        7817 => X"7C",  -- 124
        7818 => X"7B",  -- 123
        7819 => X"74",  -- 116
        7820 => X"6D",  -- 109
        7821 => X"6E",  -- 110
        7822 => X"75",  -- 117
        7823 => X"7A",  -- 122
        7824 => X"75",  -- 117
        7825 => X"66",  -- 102
        7826 => X"5C",  -- 92
        7827 => X"5C",  -- 92
        7828 => X"53",  -- 83
        7829 => X"43",  -- 67
        7830 => X"3E",  -- 62
        7831 => X"44",  -- 68
        7832 => X"40",  -- 64
        7833 => X"30",  -- 48
        7834 => X"26",  -- 38
        7835 => X"28",  -- 40
        7836 => X"2E",  -- 46
        7837 => X"2E",  -- 46
        7838 => X"2F",  -- 47
        7839 => X"33",  -- 51
        7840 => X"2A",  -- 42
        7841 => X"27",  -- 39
        7842 => X"27",  -- 39
        7843 => X"2D",  -- 45
        7844 => X"3C",  -- 60
        7845 => X"49",  -- 73
        7846 => X"49",  -- 73
        7847 => X"42",  -- 66
        7848 => X"3A",  -- 58
        7849 => X"3F",  -- 63
        7850 => X"40",  -- 64
        7851 => X"41",  -- 65
        7852 => X"4C",  -- 76
        7853 => X"5C",  -- 92
        7854 => X"60",  -- 96
        7855 => X"57",  -- 87
        7856 => X"5E",  -- 94
        7857 => X"58",  -- 88
        7858 => X"5F",  -- 95
        7859 => X"72",  -- 114
        7860 => X"79",  -- 121
        7861 => X"70",  -- 112
        7862 => X"6A",  -- 106
        7863 => X"6E",  -- 110
        7864 => X"6A",  -- 106
        7865 => X"6F",  -- 111
        7866 => X"73",  -- 115
        7867 => X"75",  -- 117
        7868 => X"75",  -- 117
        7869 => X"77",  -- 119
        7870 => X"7C",  -- 124
        7871 => X"80",  -- 128
        7872 => X"7F",  -- 127
        7873 => X"7D",  -- 125
        7874 => X"7A",  -- 122
        7875 => X"78",  -- 120
        7876 => X"77",  -- 119
        7877 => X"7A",  -- 122
        7878 => X"7E",  -- 126
        7879 => X"81",  -- 129
        7880 => X"81",  -- 129
        7881 => X"85",  -- 133
        7882 => X"8F",  -- 143
        7883 => X"96",  -- 150
        7884 => X"95",  -- 149
        7885 => X"90",  -- 144
        7886 => X"91",  -- 145
        7887 => X"96",  -- 150
        7888 => X"93",  -- 147
        7889 => X"96",  -- 150
        7890 => X"98",  -- 152
        7891 => X"9A",  -- 154
        7892 => X"A2",  -- 162
        7893 => X"AF",  -- 175
        7894 => X"B2",  -- 178
        7895 => X"AE",  -- 174
        7896 => X"B6",  -- 182
        7897 => X"B8",  -- 184
        7898 => X"BB",  -- 187
        7899 => X"BD",  -- 189
        7900 => X"BD",  -- 189
        7901 => X"BB",  -- 187
        7902 => X"B9",  -- 185
        7903 => X"B8",  -- 184
        7904 => X"AF",  -- 175
        7905 => X"A9",  -- 169
        7906 => X"9A",  -- 154
        7907 => X"89",  -- 137
        7908 => X"87",  -- 135
        7909 => X"8D",  -- 141
        7910 => X"91",  -- 145
        7911 => X"8D",  -- 141
        7912 => X"8F",  -- 143
        7913 => X"88",  -- 136
        7914 => X"87",  -- 135
        7915 => X"92",  -- 146
        7916 => X"98",  -- 152
        7917 => X"95",  -- 149
        7918 => X"95",  -- 149
        7919 => X"99",  -- 153
        7920 => X"A5",  -- 165
        7921 => X"AA",  -- 170
        7922 => X"AB",  -- 171
        7923 => X"A8",  -- 168
        7924 => X"A8",  -- 168
        7925 => X"AB",  -- 171
        7926 => X"AA",  -- 170
        7927 => X"A7",  -- 167
        7928 => X"A5",  -- 165
        7929 => X"A8",  -- 168
        7930 => X"AD",  -- 173
        7931 => X"B1",  -- 177
        7932 => X"B3",  -- 179
        7933 => X"B2",  -- 178
        7934 => X"B1",  -- 177
        7935 => X"AF",  -- 175
        7936 => X"A7",  -- 167
        7937 => X"AF",  -- 175
        7938 => X"B7",  -- 183
        7939 => X"B9",  -- 185
        7940 => X"B7",  -- 183
        7941 => X"B7",  -- 183
        7942 => X"B3",  -- 179
        7943 => X"AF",  -- 175
        7944 => X"A5",  -- 165
        7945 => X"98",  -- 152
        7946 => X"8C",  -- 140
        7947 => X"7A",  -- 122
        7948 => X"5D",  -- 93
        7949 => X"4C",  -- 76
        7950 => X"62",  -- 98
        7951 => X"85",  -- 133
        7952 => X"87",  -- 135
        7953 => X"8D",  -- 141
        7954 => X"9B",  -- 155
        7955 => X"A7",  -- 167
        7956 => X"A8",  -- 168
        7957 => X"A0",  -- 160
        7958 => X"9E",  -- 158
        7959 => X"A4",  -- 164
        7960 => X"A0",  -- 160
        7961 => X"9F",  -- 159
        7962 => X"9F",  -- 159
        7963 => X"9F",  -- 159
        7964 => X"9F",  -- 159
        7965 => X"9D",  -- 157
        7966 => X"9A",  -- 154
        7967 => X"98",  -- 152
        7968 => X"8F",  -- 143
        7969 => X"87",  -- 135
        7970 => X"7D",  -- 125
        7971 => X"74",  -- 116
        7972 => X"6F",  -- 111
        7973 => X"68",  -- 104
        7974 => X"5E",  -- 94
        7975 => X"56",  -- 86
        7976 => X"52",  -- 82
        7977 => X"63",  -- 99
        7978 => X"7C",  -- 124
        7979 => X"97",  -- 151
        7980 => X"AC",  -- 172
        7981 => X"B4",  -- 180
        7982 => X"B4",  -- 180
        7983 => X"B1",  -- 177
        7984 => X"B5",  -- 181
        7985 => X"B8",  -- 184
        7986 => X"BB",  -- 187
        7987 => X"B9",  -- 185
        7988 => X"B5",  -- 181
        7989 => X"B4",  -- 180
        7990 => X"B4",  -- 180
        7991 => X"B5",  -- 181
        7992 => X"BC",  -- 188
        7993 => X"BB",  -- 187
        7994 => X"C3",  -- 195
        7995 => X"BB",  -- 187
        7996 => X"A1",  -- 161
        7997 => X"9E",  -- 158
        7998 => X"AD",  -- 173
        7999 => X"AD",  -- 173
        8000 => X"3D",  -- 61
        8001 => X"3C",  -- 60
        8002 => X"3C",  -- 60
        8003 => X"3C",  -- 60
        8004 => X"3D",  -- 61
        8005 => X"3D",  -- 61
        8006 => X"3E",  -- 62
        8007 => X"3F",  -- 63
        8008 => X"3E",  -- 62
        8009 => X"3E",  -- 62
        8010 => X"3F",  -- 63
        8011 => X"3F",  -- 63
        8012 => X"3F",  -- 63
        8013 => X"3F",  -- 63
        8014 => X"3E",  -- 62
        8015 => X"3E",  -- 62
        8016 => X"3E",  -- 62
        8017 => X"3E",  -- 62
        8018 => X"3E",  -- 62
        8019 => X"3E",  -- 62
        8020 => X"3E",  -- 62
        8021 => X"3D",  -- 61
        8022 => X"3D",  -- 61
        8023 => X"3D",  -- 61
        8024 => X"3E",  -- 62
        8025 => X"3E",  -- 62
        8026 => X"3E",  -- 62
        8027 => X"3E",  -- 62
        8028 => X"3E",  -- 62
        8029 => X"3D",  -- 61
        8030 => X"3D",  -- 61
        8031 => X"3D",  -- 61
        8032 => X"3C",  -- 60
        8033 => X"3C",  -- 60
        8034 => X"3C",  -- 60
        8035 => X"3B",  -- 59
        8036 => X"3A",  -- 58
        8037 => X"37",  -- 55
        8038 => X"35",  -- 53
        8039 => X"34",  -- 52
        8040 => X"34",  -- 52
        8041 => X"33",  -- 51
        8042 => X"33",  -- 51
        8043 => X"33",  -- 51
        8044 => X"34",  -- 52
        8045 => X"34",  -- 52
        8046 => X"34",  -- 52
        8047 => X"34",  -- 52
        8048 => X"34",  -- 52
        8049 => X"33",  -- 51
        8050 => X"31",  -- 49
        8051 => X"2E",  -- 46
        8052 => X"30",  -- 48
        8053 => X"34",  -- 52
        8054 => X"3B",  -- 59
        8055 => X"3F",  -- 63
        8056 => X"49",  -- 73
        8057 => X"52",  -- 82
        8058 => X"5C",  -- 92
        8059 => X"66",  -- 102
        8060 => X"69",  -- 105
        8061 => X"6D",  -- 109
        8062 => X"72",  -- 114
        8063 => X"76",  -- 118
        8064 => X"7B",  -- 123
        8065 => X"7E",  -- 126
        8066 => X"81",  -- 129
        8067 => X"84",  -- 132
        8068 => X"85",  -- 133
        8069 => X"84",  -- 132
        8070 => X"81",  -- 129
        8071 => X"7E",  -- 126
        8072 => X"76",  -- 118
        8073 => X"7A",  -- 122
        8074 => X"79",  -- 121
        8075 => X"7D",  -- 125
        8076 => X"8F",  -- 143
        8077 => X"9E",  -- 158
        8078 => X"A1",  -- 161
        8079 => X"A3",  -- 163
        8080 => X"A4",  -- 164
        8081 => X"A1",  -- 161
        8082 => X"A4",  -- 164
        8083 => X"97",  -- 151
        8084 => X"A0",  -- 160
        8085 => X"9A",  -- 154
        8086 => X"9F",  -- 159
        8087 => X"96",  -- 150
        8088 => X"96",  -- 150
        8089 => X"8C",  -- 140
        8090 => X"93",  -- 147
        8091 => X"91",  -- 145
        8092 => X"9E",  -- 158
        8093 => X"91",  -- 145
        8094 => X"94",  -- 148
        8095 => X"92",  -- 146
        8096 => X"94",  -- 148
        8097 => X"9B",  -- 155
        8098 => X"98",  -- 152
        8099 => X"9C",  -- 156
        8100 => X"9A",  -- 154
        8101 => X"99",  -- 153
        8102 => X"A1",  -- 161
        8103 => X"97",  -- 151
        8104 => X"90",  -- 144
        8105 => X"7A",  -- 122
        8106 => X"78",  -- 120
        8107 => X"82",  -- 130
        8108 => X"86",  -- 134
        8109 => X"92",  -- 146
        8110 => X"8B",  -- 139
        8111 => X"8B",  -- 139
        8112 => X"94",  -- 148
        8113 => X"99",  -- 153
        8114 => X"94",  -- 148
        8115 => X"92",  -- 146
        8116 => X"7B",  -- 123
        8117 => X"70",  -- 112
        8118 => X"90",  -- 144
        8119 => X"7E",  -- 126
        8120 => X"81",  -- 129
        8121 => X"92",  -- 146
        8122 => X"8D",  -- 141
        8123 => X"92",  -- 146
        8124 => X"94",  -- 148
        8125 => X"86",  -- 134
        8126 => X"7E",  -- 126
        8127 => X"75",  -- 117
        8128 => X"72",  -- 114
        8129 => X"77",  -- 119
        8130 => X"74",  -- 116
        8131 => X"71",  -- 113
        8132 => X"77",  -- 119
        8133 => X"78",  -- 120
        8134 => X"75",  -- 117
        8135 => X"79",  -- 121
        8136 => X"7C",  -- 124
        8137 => X"80",  -- 128
        8138 => X"80",  -- 128
        8139 => X"7B",  -- 123
        8140 => X"77",  -- 119
        8141 => X"7A",  -- 122
        8142 => X"80",  -- 128
        8143 => X"83",  -- 131
        8144 => X"77",  -- 119
        8145 => X"6F",  -- 111
        8146 => X"6B",  -- 107
        8147 => X"6A",  -- 106
        8148 => X"65",  -- 101
        8149 => X"5D",  -- 93
        8150 => X"58",  -- 88
        8151 => X"5A",  -- 90
        8152 => X"3A",  -- 58
        8153 => X"36",  -- 54
        8154 => X"34",  -- 52
        8155 => X"32",  -- 50
        8156 => X"2F",  -- 47
        8157 => X"2B",  -- 43
        8158 => X"2C",  -- 44
        8159 => X"2F",  -- 47
        8160 => X"2A",  -- 42
        8161 => X"31",  -- 49
        8162 => X"34",  -- 52
        8163 => X"30",  -- 48
        8164 => X"2C",  -- 44
        8165 => X"31",  -- 49
        8166 => X"39",  -- 57
        8167 => X"3E",  -- 62
        8168 => X"3B",  -- 59
        8169 => X"41",  -- 65
        8170 => X"4A",  -- 74
        8171 => X"50",  -- 80
        8172 => X"54",  -- 84
        8173 => X"54",  -- 84
        8174 => X"55",  -- 85
        8175 => X"58",  -- 88
        8176 => X"5E",  -- 94
        8177 => X"63",  -- 99
        8178 => X"6A",  -- 106
        8179 => X"6C",  -- 108
        8180 => X"69",  -- 105
        8181 => X"66",  -- 102
        8182 => X"6B",  -- 107
        8183 => X"71",  -- 113
        8184 => X"6C",  -- 108
        8185 => X"6F",  -- 111
        8186 => X"72",  -- 114
        8187 => X"73",  -- 115
        8188 => X"72",  -- 114
        8189 => X"74",  -- 116
        8190 => X"79",  -- 121
        8191 => X"7D",  -- 125
        8192 => X"78",  -- 120
        8193 => X"78",  -- 120
        8194 => X"76",  -- 118
        8195 => X"73",  -- 115
        8196 => X"73",  -- 115
        8197 => X"77",  -- 119
        8198 => X"7D",  -- 125
        8199 => X"83",  -- 131
        8200 => X"7A",  -- 122
        8201 => X"7F",  -- 127
        8202 => X"88",  -- 136
        8203 => X"90",  -- 144
        8204 => X"91",  -- 145
        8205 => X"8E",  -- 142
        8206 => X"91",  -- 145
        8207 => X"97",  -- 151
        8208 => X"92",  -- 146
        8209 => X"98",  -- 152
        8210 => X"9B",  -- 155
        8211 => X"9D",  -- 157
        8212 => X"A2",  -- 162
        8213 => X"AA",  -- 170
        8214 => X"B0",  -- 176
        8215 => X"B2",  -- 178
        8216 => X"B2",  -- 178
        8217 => X"B5",  -- 181
        8218 => X"B8",  -- 184
        8219 => X"B9",  -- 185
        8220 => X"B9",  -- 185
        8221 => X"B8",  -- 184
        8222 => X"B7",  -- 183
        8223 => X"B6",  -- 182
        8224 => X"B6",  -- 182
        8225 => X"B0",  -- 176
        8226 => X"A4",  -- 164
        8227 => X"97",  -- 151
        8228 => X"92",  -- 146
        8229 => X"94",  -- 148
        8230 => X"94",  -- 148
        8231 => X"93",  -- 147
        8232 => X"90",  -- 144
        8233 => X"8D",  -- 141
        8234 => X"90",  -- 144
        8235 => X"98",  -- 152
        8236 => X"98",  -- 152
        8237 => X"94",  -- 148
        8238 => X"97",  -- 151
        8239 => X"9F",  -- 159
        8240 => X"AB",  -- 171
        8241 => X"AD",  -- 173
        8242 => X"AD",  -- 173
        8243 => X"AA",  -- 170
        8244 => X"A9",  -- 169
        8245 => X"AA",  -- 170
        8246 => X"A7",  -- 167
        8247 => X"A2",  -- 162
        8248 => X"A7",  -- 167
        8249 => X"A9",  -- 169
        8250 => X"AD",  -- 173
        8251 => X"B0",  -- 176
        8252 => X"B1",  -- 177
        8253 => X"B0",  -- 176
        8254 => X"AD",  -- 173
        8255 => X"AA",  -- 170
        8256 => X"AD",  -- 173
        8257 => X"B0",  -- 176
        8258 => X"B2",  -- 178
        8259 => X"B0",  -- 176
        8260 => X"AF",  -- 175
        8261 => X"B1",  -- 177
        8262 => X"AD",  -- 173
        8263 => X"AB",  -- 171
        8264 => X"A3",  -- 163
        8265 => X"9E",  -- 158
        8266 => X"96",  -- 150
        8267 => X"88",  -- 136
        8268 => X"6E",  -- 110
        8269 => X"57",  -- 87
        8270 => X"5C",  -- 92
        8271 => X"6D",  -- 109
        8272 => X"6C",  -- 108
        8273 => X"76",  -- 118
        8274 => X"88",  -- 136
        8275 => X"97",  -- 151
        8276 => X"9D",  -- 157
        8277 => X"9E",  -- 158
        8278 => X"A2",  -- 162
        8279 => X"A7",  -- 167
        8280 => X"A1",  -- 161
        8281 => X"9F",  -- 159
        8282 => X"9C",  -- 156
        8283 => X"9C",  -- 156
        8284 => X"9C",  -- 156
        8285 => X"9F",  -- 159
        8286 => X"A1",  -- 161
        8287 => X"A3",  -- 163
        8288 => X"95",  -- 149
        8289 => X"8C",  -- 140
        8290 => X"83",  -- 131
        8291 => X"7D",  -- 125
        8292 => X"78",  -- 120
        8293 => X"6E",  -- 110
        8294 => X"5D",  -- 93
        8295 => X"50",  -- 80
        8296 => X"50",  -- 80
        8297 => X"5C",  -- 92
        8298 => X"70",  -- 112
        8299 => X"8C",  -- 140
        8300 => X"A6",  -- 166
        8301 => X"B4",  -- 180
        8302 => X"B4",  -- 180
        8303 => X"B0",  -- 176
        8304 => X"BA",  -- 186
        8305 => X"BB",  -- 187
        8306 => X"BA",  -- 186
        8307 => X"B6",  -- 182
        8308 => X"B1",  -- 177
        8309 => X"B0",  -- 176
        8310 => X"B2",  -- 178
        8311 => X"B4",  -- 180
        8312 => X"BE",  -- 190
        8313 => X"BA",  -- 186
        8314 => X"BD",  -- 189
        8315 => X"B0",  -- 176
        8316 => X"99",  -- 153
        8317 => X"9B",  -- 155
        8318 => X"AE",  -- 174
        8319 => X"B1",  -- 177
        8320 => X"3C",  -- 60
        8321 => X"3C",  -- 60
        8322 => X"3C",  -- 60
        8323 => X"3C",  -- 60
        8324 => X"3D",  -- 61
        8325 => X"3E",  -- 62
        8326 => X"3E",  -- 62
        8327 => X"3F",  -- 63
        8328 => X"3E",  -- 62
        8329 => X"3F",  -- 63
        8330 => X"3F",  -- 63
        8331 => X"40",  -- 64
        8332 => X"40",  -- 64
        8333 => X"3F",  -- 63
        8334 => X"3F",  -- 63
        8335 => X"3E",  -- 62
        8336 => X"3F",  -- 63
        8337 => X"3F",  -- 63
        8338 => X"3E",  -- 62
        8339 => X"3E",  -- 62
        8340 => X"3E",  -- 62
        8341 => X"3E",  -- 62
        8342 => X"3D",  -- 61
        8343 => X"3D",  -- 61
        8344 => X"3E",  -- 62
        8345 => X"3E",  -- 62
        8346 => X"3E",  -- 62
        8347 => X"3E",  -- 62
        8348 => X"3D",  -- 61
        8349 => X"3D",  -- 61
        8350 => X"3D",  -- 61
        8351 => X"3D",  -- 61
        8352 => X"3C",  -- 60
        8353 => X"3C",  -- 60
        8354 => X"3C",  -- 60
        8355 => X"3B",  -- 59
        8356 => X"3A",  -- 58
        8357 => X"38",  -- 56
        8358 => X"36",  -- 54
        8359 => X"35",  -- 53
        8360 => X"35",  -- 53
        8361 => X"34",  -- 52
        8362 => X"33",  -- 51
        8363 => X"33",  -- 51
        8364 => X"33",  -- 51
        8365 => X"32",  -- 50
        8366 => X"33",  -- 51
        8367 => X"32",  -- 50
        8368 => X"32",  -- 50
        8369 => X"31",  -- 49
        8370 => X"30",  -- 48
        8371 => X"32",  -- 50
        8372 => X"39",  -- 57
        8373 => X"44",  -- 68
        8374 => X"50",  -- 80
        8375 => X"59",  -- 89
        8376 => X"62",  -- 98
        8377 => X"68",  -- 104
        8378 => X"71",  -- 113
        8379 => X"78",  -- 120
        8380 => X"7D",  -- 125
        8381 => X"81",  -- 129
        8382 => X"85",  -- 133
        8383 => X"86",  -- 134
        8384 => X"8B",  -- 139
        8385 => X"8B",  -- 139
        8386 => X"8D",  -- 141
        8387 => X"8E",  -- 142
        8388 => X"8B",  -- 139
        8389 => X"88",  -- 136
        8390 => X"81",  -- 129
        8391 => X"7D",  -- 125
        8392 => X"77",  -- 119
        8393 => X"77",  -- 119
        8394 => X"76",  -- 118
        8395 => X"7A",  -- 122
        8396 => X"90",  -- 144
        8397 => X"A5",  -- 165
        8398 => X"A6",  -- 166
        8399 => X"9C",  -- 156
        8400 => X"A0",  -- 160
        8401 => X"9B",  -- 155
        8402 => X"9C",  -- 156
        8403 => X"90",  -- 144
        8404 => X"94",  -- 148
        8405 => X"8C",  -- 140
        8406 => X"8C",  -- 140
        8407 => X"84",  -- 132
        8408 => X"7E",  -- 126
        8409 => X"7E",  -- 126
        8410 => X"84",  -- 132
        8411 => X"7E",  -- 126
        8412 => X"84",  -- 132
        8413 => X"83",  -- 131
        8414 => X"91",  -- 145
        8415 => X"94",  -- 148
        8416 => X"93",  -- 147
        8417 => X"98",  -- 152
        8418 => X"91",  -- 145
        8419 => X"96",  -- 150
        8420 => X"96",  -- 150
        8421 => X"92",  -- 146
        8422 => X"96",  -- 150
        8423 => X"8B",  -- 139
        8424 => X"8D",  -- 141
        8425 => X"79",  -- 121
        8426 => X"83",  -- 131
        8427 => X"84",  -- 132
        8428 => X"8C",  -- 140
        8429 => X"8C",  -- 140
        8430 => X"8A",  -- 138
        8431 => X"8B",  -- 139
        8432 => X"97",  -- 151
        8433 => X"99",  -- 153
        8434 => X"82",  -- 130
        8435 => X"79",  -- 121
        8436 => X"5B",  -- 91
        8437 => X"5F",  -- 95
        8438 => X"7D",  -- 125
        8439 => X"73",  -- 115
        8440 => X"72",  -- 114
        8441 => X"87",  -- 135
        8442 => X"86",  -- 134
        8443 => X"89",  -- 137
        8444 => X"8B",  -- 139
        8445 => X"82",  -- 130
        8446 => X"7F",  -- 127
        8447 => X"78",  -- 120
        8448 => X"72",  -- 114
        8449 => X"7B",  -- 123
        8450 => X"78",  -- 120
        8451 => X"70",  -- 112
        8452 => X"77",  -- 119
        8453 => X"80",  -- 128
        8454 => X"7E",  -- 126
        8455 => X"7B",  -- 123
        8456 => X"7E",  -- 126
        8457 => X"81",  -- 129
        8458 => X"82",  -- 130
        8459 => X"7F",  -- 127
        8460 => X"7D",  -- 125
        8461 => X"80",  -- 128
        8462 => X"81",  -- 129
        8463 => X"80",  -- 128
        8464 => X"7F",  -- 127
        8465 => X"7E",  -- 126
        8466 => X"7B",  -- 123
        8467 => X"77",  -- 119
        8468 => X"70",  -- 112
        8469 => X"6A",  -- 106
        8470 => X"63",  -- 99
        8471 => X"5D",  -- 93
        8472 => X"46",  -- 70
        8473 => X"4C",  -- 76
        8474 => X"4B",  -- 75
        8475 => X"42",  -- 66
        8476 => X"38",  -- 56
        8477 => X"35",  -- 53
        8478 => X"3A",  -- 58
        8479 => X"3D",  -- 61
        8480 => X"39",  -- 57
        8481 => X"39",  -- 57
        8482 => X"37",  -- 55
        8483 => X"33",  -- 51
        8484 => X"32",  -- 50
        8485 => X"36",  -- 54
        8486 => X"35",  -- 53
        8487 => X"33",  -- 51
        8488 => X"3A",  -- 58
        8489 => X"39",  -- 57
        8490 => X"44",  -- 68
        8491 => X"55",  -- 85
        8492 => X"5A",  -- 90
        8493 => X"55",  -- 85
        8494 => X"57",  -- 87
        8495 => X"60",  -- 96
        8496 => X"61",  -- 97
        8497 => X"6B",  -- 107
        8498 => X"70",  -- 112
        8499 => X"69",  -- 105
        8500 => X"64",  -- 100
        8501 => X"67",  -- 103
        8502 => X"6B",  -- 107
        8503 => X"6B",  -- 107
        8504 => X"66",  -- 102
        8505 => X"68",  -- 104
        8506 => X"6A",  -- 106
        8507 => X"6B",  -- 107
        8508 => X"6B",  -- 107
        8509 => X"6D",  -- 109
        8510 => X"72",  -- 114
        8511 => X"77",  -- 119
        8512 => X"74",  -- 116
        8513 => X"74",  -- 116
        8514 => X"74",  -- 116
        8515 => X"71",  -- 113
        8516 => X"70",  -- 112
        8517 => X"73",  -- 115
        8518 => X"7A",  -- 122
        8519 => X"81",  -- 129
        8520 => X"7D",  -- 125
        8521 => X"81",  -- 129
        8522 => X"88",  -- 136
        8523 => X"8D",  -- 141
        8524 => X"8C",  -- 140
        8525 => X"89",  -- 137
        8526 => X"8B",  -- 139
        8527 => X"8F",  -- 143
        8528 => X"92",  -- 146
        8529 => X"96",  -- 150
        8530 => X"9C",  -- 156
        8531 => X"A2",  -- 162
        8532 => X"A2",  -- 162
        8533 => X"A4",  -- 164
        8534 => X"AC",  -- 172
        8535 => X"B5",  -- 181
        8536 => X"AE",  -- 174
        8537 => X"B0",  -- 176
        8538 => X"B3",  -- 179
        8539 => X"B3",  -- 179
        8540 => X"B3",  -- 179
        8541 => X"B3",  -- 179
        8542 => X"B5",  -- 181
        8543 => X"B5",  -- 181
        8544 => X"BA",  -- 186
        8545 => X"B5",  -- 181
        8546 => X"AC",  -- 172
        8547 => X"A5",  -- 165
        8548 => X"9D",  -- 157
        8549 => X"98",  -- 152
        8550 => X"96",  -- 150
        8551 => X"99",  -- 153
        8552 => X"93",  -- 147
        8553 => X"96",  -- 150
        8554 => X"9D",  -- 157
        8555 => X"A1",  -- 161
        8556 => X"9B",  -- 155
        8557 => X"96",  -- 150
        8558 => X"9C",  -- 156
        8559 => X"A7",  -- 167
        8560 => X"AE",  -- 174
        8561 => X"AE",  -- 174
        8562 => X"AB",  -- 171
        8563 => X"A8",  -- 168
        8564 => X"A8",  -- 168
        8565 => X"A7",  -- 167
        8566 => X"A2",  -- 162
        8567 => X"9C",  -- 156
        8568 => X"A5",  -- 165
        8569 => X"A6",  -- 166
        8570 => X"AA",  -- 170
        8571 => X"AD",  -- 173
        8572 => X"B0",  -- 176
        8573 => X"AE",  -- 174
        8574 => X"AB",  -- 171
        8575 => X"A8",  -- 168
        8576 => X"B1",  -- 177
        8577 => X"B1",  -- 177
        8578 => X"AE",  -- 174
        8579 => X"AB",  -- 171
        8580 => X"AE",  -- 174
        8581 => X"B1",  -- 177
        8582 => X"B2",  -- 178
        8583 => X"B0",  -- 176
        8584 => X"A5",  -- 165
        8585 => X"A3",  -- 163
        8586 => X"9F",  -- 159
        8587 => X"94",  -- 148
        8588 => X"7F",  -- 127
        8589 => X"64",  -- 100
        8590 => X"51",  -- 81
        8591 => X"49",  -- 73
        8592 => X"51",  -- 81
        8593 => X"61",  -- 97
        8594 => X"74",  -- 116
        8595 => X"83",  -- 131
        8596 => X"8F",  -- 143
        8597 => X"9A",  -- 154
        8598 => X"A2",  -- 162
        8599 => X"A5",  -- 165
        8600 => X"9F",  -- 159
        8601 => X"9C",  -- 156
        8602 => X"99",  -- 153
        8603 => X"99",  -- 153
        8604 => X"9A",  -- 154
        8605 => X"9D",  -- 157
        8606 => X"A0",  -- 160
        8607 => X"A1",  -- 161
        8608 => X"9C",  -- 156
        8609 => X"94",  -- 148
        8610 => X"8C",  -- 140
        8611 => X"8A",  -- 138
        8612 => X"86",  -- 134
        8613 => X"7A",  -- 122
        8614 => X"62",  -- 98
        8615 => X"4F",  -- 79
        8616 => X"4C",  -- 76
        8617 => X"52",  -- 82
        8618 => X"63",  -- 99
        8619 => X"82",  -- 130
        8620 => X"A2",  -- 162
        8621 => X"B5",  -- 181
        8622 => X"B7",  -- 183
        8623 => X"B6",  -- 182
        8624 => X"BA",  -- 186
        8625 => X"BB",  -- 187
        8626 => X"BA",  -- 186
        8627 => X"B6",  -- 182
        8628 => X"B1",  -- 177
        8629 => X"AE",  -- 174
        8630 => X"AE",  -- 174
        8631 => X"AE",  -- 174
        8632 => X"BA",  -- 186
        8633 => X"B7",  -- 183
        8634 => X"B7",  -- 183
        8635 => X"A9",  -- 169
        8636 => X"97",  -- 151
        8637 => X"9C",  -- 156
        8638 => X"AD",  -- 173
        8639 => X"B1",  -- 177
        8640 => X"3C",  -- 60
        8641 => X"3C",  -- 60
        8642 => X"3C",  -- 60
        8643 => X"3C",  -- 60
        8644 => X"3D",  -- 61
        8645 => X"3E",  -- 62
        8646 => X"3F",  -- 63
        8647 => X"3F",  -- 63
        8648 => X"3F",  -- 63
        8649 => X"3F",  -- 63
        8650 => X"40",  -- 64
        8651 => X"40",  -- 64
        8652 => X"40",  -- 64
        8653 => X"40",  -- 64
        8654 => X"3F",  -- 63
        8655 => X"3F",  -- 63
        8656 => X"3F",  -- 63
        8657 => X"3F",  -- 63
        8658 => X"3F",  -- 63
        8659 => X"3E",  -- 62
        8660 => X"3E",  -- 62
        8661 => X"3E",  -- 62
        8662 => X"3E",  -- 62
        8663 => X"3E",  -- 62
        8664 => X"3E",  -- 62
        8665 => X"3E",  -- 62
        8666 => X"3E",  -- 62
        8667 => X"3D",  -- 61
        8668 => X"3D",  -- 61
        8669 => X"3D",  -- 61
        8670 => X"3D",  -- 61
        8671 => X"3C",  -- 60
        8672 => X"3A",  -- 58
        8673 => X"3A",  -- 58
        8674 => X"3B",  -- 59
        8675 => X"3B",  -- 59
        8676 => X"3B",  -- 59
        8677 => X"39",  -- 57
        8678 => X"39",  -- 57
        8679 => X"39",  -- 57
        8680 => X"38",  -- 56
        8681 => X"37",  -- 55
        8682 => X"35",  -- 53
        8683 => X"32",  -- 50
        8684 => X"30",  -- 48
        8685 => X"32",  -- 50
        8686 => X"33",  -- 51
        8687 => X"34",  -- 52
        8688 => X"36",  -- 54
        8689 => X"37",  -- 55
        8690 => X"3C",  -- 60
        8691 => X"43",  -- 67
        8692 => X"4B",  -- 75
        8693 => X"59",  -- 89
        8694 => X"65",  -- 101
        8695 => X"6E",  -- 110
        8696 => X"74",  -- 116
        8697 => X"75",  -- 117
        8698 => X"75",  -- 117
        8699 => X"78",  -- 120
        8700 => X"7D",  -- 125
        8701 => X"83",  -- 131
        8702 => X"89",  -- 137
        8703 => X"8C",  -- 140
        8704 => X"90",  -- 144
        8705 => X"8F",  -- 143
        8706 => X"8D",  -- 141
        8707 => X"8B",  -- 139
        8708 => X"8A",  -- 138
        8709 => X"87",  -- 135
        8710 => X"83",  -- 131
        8711 => X"7F",  -- 127
        8712 => X"84",  -- 132
        8713 => X"7F",  -- 127
        8714 => X"7D",  -- 125
        8715 => X"7F",  -- 127
        8716 => X"8E",  -- 142
        8717 => X"9F",  -- 159
        8718 => X"A0",  -- 160
        8719 => X"91",  -- 145
        8720 => X"90",  -- 144
        8721 => X"87",  -- 135
        8722 => X"83",  -- 131
        8723 => X"76",  -- 118
        8724 => X"7C",  -- 124
        8725 => X"71",  -- 113
        8726 => X"6F",  -- 111
        8727 => X"66",  -- 102
        8728 => X"5B",  -- 91
        8729 => X"61",  -- 97
        8730 => X"63",  -- 99
        8731 => X"5E",  -- 94
        8732 => X"65",  -- 101
        8733 => X"73",  -- 115
        8734 => X"85",  -- 133
        8735 => X"8D",  -- 141
        8736 => X"8A",  -- 138
        8737 => X"90",  -- 144
        8738 => X"87",  -- 135
        8739 => X"8C",  -- 140
        8740 => X"91",  -- 145
        8741 => X"8A",  -- 138
        8742 => X"8B",  -- 139
        8743 => X"84",  -- 132
        8744 => X"86",  -- 134
        8745 => X"72",  -- 114
        8746 => X"82",  -- 130
        8747 => X"7E",  -- 126
        8748 => X"88",  -- 136
        8749 => X"80",  -- 128
        8750 => X"7F",  -- 127
        8751 => X"7B",  -- 123
        8752 => X"8E",  -- 142
        8753 => X"86",  -- 134
        8754 => X"5C",  -- 92
        8755 => X"4F",  -- 79
        8756 => X"39",  -- 57
        8757 => X"4E",  -- 78
        8758 => X"62",  -- 98
        8759 => X"5B",  -- 91
        8760 => X"64",  -- 100
        8761 => X"77",  -- 119
        8762 => X"75",  -- 117
        8763 => X"78",  -- 120
        8764 => X"7D",  -- 125
        8765 => X"7D",  -- 125
        8766 => X"84",  -- 132
        8767 => X"82",  -- 130
        8768 => X"79",  -- 121
        8769 => X"80",  -- 128
        8770 => X"7B",  -- 123
        8771 => X"76",  -- 118
        8772 => X"7D",  -- 125
        8773 => X"80",  -- 128
        8774 => X"7C",  -- 124
        8775 => X"7B",  -- 123
        8776 => X"7E",  -- 126
        8777 => X"81",  -- 129
        8778 => X"81",  -- 129
        8779 => X"80",  -- 128
        8780 => X"80",  -- 128
        8781 => X"82",  -- 130
        8782 => X"80",  -- 128
        8783 => X"7B",  -- 123
        8784 => X"84",  -- 132
        8785 => X"86",  -- 134
        8786 => X"82",  -- 130
        8787 => X"79",  -- 121
        8788 => X"74",  -- 116
        8789 => X"70",  -- 112
        8790 => X"69",  -- 105
        8791 => X"5F",  -- 95
        8792 => X"5E",  -- 94
        8793 => X"60",  -- 96
        8794 => X"5A",  -- 90
        8795 => X"4C",  -- 76
        8796 => X"45",  -- 69
        8797 => X"4D",  -- 77
        8798 => X"56",  -- 86
        8799 => X"5A",  -- 90
        8800 => X"51",  -- 81
        8801 => X"4A",  -- 74
        8802 => X"40",  -- 64
        8803 => X"3C",  -- 60
        8804 => X"3C",  -- 60
        8805 => X"3E",  -- 62
        8806 => X"35",  -- 53
        8807 => X"2A",  -- 42
        8808 => X"3A",  -- 58
        8809 => X"36",  -- 54
        8810 => X"3B",  -- 59
        8811 => X"4B",  -- 75
        8812 => X"58",  -- 88
        8813 => X"5B",  -- 91
        8814 => X"5E",  -- 94
        8815 => X"64",  -- 100
        8816 => X"64",  -- 100
        8817 => X"66",  -- 102
        8818 => X"69",  -- 105
        8819 => X"6B",  -- 107
        8820 => X"6E",  -- 110
        8821 => X"6F",  -- 111
        8822 => X"68",  -- 104
        8823 => X"5F",  -- 95
        8824 => X"64",  -- 100
        8825 => X"65",  -- 101
        8826 => X"66",  -- 102
        8827 => X"67",  -- 103
        8828 => X"68",  -- 104
        8829 => X"6B",  -- 107
        8830 => X"70",  -- 112
        8831 => X"74",  -- 116
        8832 => X"73",  -- 115
        8833 => X"75",  -- 117
        8834 => X"77",  -- 119
        8835 => X"74",  -- 116
        8836 => X"71",  -- 113
        8837 => X"71",  -- 113
        8838 => X"76",  -- 118
        8839 => X"7B",  -- 123
        8840 => X"7C",  -- 124
        8841 => X"80",  -- 128
        8842 => X"85",  -- 133
        8843 => X"88",  -- 136
        8844 => X"87",  -- 135
        8845 => X"87",  -- 135
        8846 => X"87",  -- 135
        8847 => X"89",  -- 137
        8848 => X"92",  -- 146
        8849 => X"92",  -- 146
        8850 => X"99",  -- 153
        8851 => X"A2",  -- 162
        8852 => X"A4",  -- 164
        8853 => X"A0",  -- 160
        8854 => X"A5",  -- 165
        8855 => X"AF",  -- 175
        8856 => X"AC",  -- 172
        8857 => X"AE",  -- 174
        8858 => X"B0",  -- 176
        8859 => X"B1",  -- 177
        8860 => X"B0",  -- 176
        8861 => X"B2",  -- 178
        8862 => X"B5",  -- 181
        8863 => X"B6",  -- 182
        8864 => X"B8",  -- 184
        8865 => X"B2",  -- 178
        8866 => X"AD",  -- 173
        8867 => X"AA",  -- 170
        8868 => X"A2",  -- 162
        8869 => X"98",  -- 152
        8870 => X"98",  -- 152
        8871 => X"9F",  -- 159
        8872 => X"9B",  -- 155
        8873 => X"9F",  -- 159
        8874 => X"A5",  -- 165
        8875 => X"A7",  -- 167
        8876 => X"A1",  -- 161
        8877 => X"9C",  -- 156
        8878 => X"A2",  -- 162
        8879 => X"AD",  -- 173
        8880 => X"AB",  -- 171
        8881 => X"A9",  -- 169
        8882 => X"A6",  -- 166
        8883 => X"A5",  -- 165
        8884 => X"A5",  -- 165
        8885 => X"A4",  -- 164
        8886 => X"9F",  -- 159
        8887 => X"9A",  -- 154
        8888 => X"A0",  -- 160
        8889 => X"A2",  -- 162
        8890 => X"A5",  -- 165
        8891 => X"A9",  -- 169
        8892 => X"AE",  -- 174
        8893 => X"AE",  -- 174
        8894 => X"AC",  -- 172
        8895 => X"A9",  -- 169
        8896 => X"B0",  -- 176
        8897 => X"AF",  -- 175
        8898 => X"AC",  -- 172
        8899 => X"AB",  -- 171
        8900 => X"AF",  -- 175
        8901 => X"B3",  -- 179
        8902 => X"B1",  -- 177
        8903 => X"AC",  -- 172
        8904 => X"A1",  -- 161
        8905 => X"A5",  -- 165
        8906 => X"A2",  -- 162
        8907 => X"9A",  -- 154
        8908 => X"8D",  -- 141
        8909 => X"79",  -- 121
        8910 => X"5C",  -- 92
        8911 => X"45",  -- 69
        8912 => X"47",  -- 71
        8913 => X"58",  -- 88
        8914 => X"68",  -- 104
        8915 => X"75",  -- 117
        8916 => X"84",  -- 132
        8917 => X"96",  -- 150
        8918 => X"9F",  -- 159
        8919 => X"A0",  -- 160
        8920 => X"9E",  -- 158
        8921 => X"9F",  -- 159
        8922 => X"9E",  -- 158
        8923 => X"9F",  -- 159
        8924 => X"9F",  -- 159
        8925 => X"9E",  -- 158
        8926 => X"9B",  -- 155
        8927 => X"9A",  -- 154
        8928 => X"A3",  -- 163
        8929 => X"9D",  -- 157
        8930 => X"98",  -- 152
        8931 => X"97",  -- 151
        8932 => X"91",  -- 145
        8933 => X"7F",  -- 127
        8934 => X"67",  -- 103
        8935 => X"54",  -- 84
        8936 => X"54",  -- 84
        8937 => X"57",  -- 87
        8938 => X"67",  -- 103
        8939 => X"82",  -- 130
        8940 => X"9F",  -- 159
        8941 => X"B1",  -- 177
        8942 => X"B6",  -- 182
        8943 => X"B4",  -- 180
        8944 => X"B2",  -- 178
        8945 => X"B4",  -- 180
        8946 => X"B6",  -- 182
        8947 => X"B5",  -- 181
        8948 => X"AF",  -- 175
        8949 => X"AA",  -- 170
        8950 => X"A7",  -- 167
        8951 => X"A5",  -- 165
        8952 => X"B2",  -- 178
        8953 => X"B5",  -- 181
        8954 => X"B5",  -- 181
        8955 => X"A8",  -- 168
        8956 => X"9F",  -- 159
        8957 => X"A2",  -- 162
        8958 => X"AA",  -- 170
        8959 => X"AC",  -- 172
        8960 => X"3B",  -- 59
        8961 => X"3B",  -- 59
        8962 => X"3B",  -- 59
        8963 => X"3C",  -- 60
        8964 => X"3D",  -- 61
        8965 => X"3E",  -- 62
        8966 => X"3F",  -- 63
        8967 => X"40",  -- 64
        8968 => X"40",  -- 64
        8969 => X"40",  -- 64
        8970 => X"41",  -- 65
        8971 => X"41",  -- 65
        8972 => X"41",  -- 65
        8973 => X"41",  -- 65
        8974 => X"40",  -- 64
        8975 => X"40",  -- 64
        8976 => X"3F",  -- 63
        8977 => X"3F",  -- 63
        8978 => X"3F",  -- 63
        8979 => X"3F",  -- 63
        8980 => X"3F",  -- 63
        8981 => X"3E",  -- 62
        8982 => X"3E",  -- 62
        8983 => X"3E",  -- 62
        8984 => X"3E",  -- 62
        8985 => X"3D",  -- 61
        8986 => X"3D",  -- 61
        8987 => X"3D",  -- 61
        8988 => X"3D",  -- 61
        8989 => X"3C",  -- 60
        8990 => X"3C",  -- 60
        8991 => X"3C",  -- 60
        8992 => X"3A",  -- 58
        8993 => X"3A",  -- 58
        8994 => X"39",  -- 57
        8995 => X"39",  -- 57
        8996 => X"39",  -- 57
        8997 => X"38",  -- 56
        8998 => X"38",  -- 56
        8999 => X"39",  -- 57
        9000 => X"34",  -- 52
        9001 => X"34",  -- 52
        9002 => X"33",  -- 51
        9003 => X"31",  -- 49
        9004 => X"32",  -- 50
        9005 => X"36",  -- 54
        9006 => X"3C",  -- 60
        9007 => X"40",  -- 64
        9008 => X"44",  -- 68
        9009 => X"49",  -- 73
        9010 => X"53",  -- 83
        9011 => X"5D",  -- 93
        9012 => X"64",  -- 100
        9013 => X"6A",  -- 106
        9014 => X"6F",  -- 111
        9015 => X"73",  -- 115
        9016 => X"77",  -- 119
        9017 => X"76",  -- 118
        9018 => X"74",  -- 116
        9019 => X"75",  -- 117
        9020 => X"79",  -- 121
        9021 => X"80",  -- 128
        9022 => X"86",  -- 134
        9023 => X"8B",  -- 139
        9024 => X"8D",  -- 141
        9025 => X"8A",  -- 138
        9026 => X"87",  -- 135
        9027 => X"85",  -- 133
        9028 => X"86",  -- 134
        9029 => X"87",  -- 135
        9030 => X"88",  -- 136
        9031 => X"89",  -- 137
        9032 => X"89",  -- 137
        9033 => X"84",  -- 132
        9034 => X"89",  -- 137
        9035 => X"8A",  -- 138
        9036 => X"89",  -- 137
        9037 => X"8C",  -- 140
        9038 => X"89",  -- 137
        9039 => X"78",  -- 120
        9040 => X"70",  -- 112
        9041 => X"61",  -- 97
        9042 => X"5B",  -- 91
        9043 => X"50",  -- 80
        9044 => X"5B",  -- 91
        9045 => X"54",  -- 84
        9046 => X"55",  -- 85
        9047 => X"4C",  -- 76
        9048 => X"3D",  -- 61
        9049 => X"43",  -- 67
        9050 => X"42",  -- 66
        9051 => X"40",  -- 64
        9052 => X"4A",  -- 74
        9053 => X"63",  -- 99
        9054 => X"73",  -- 115
        9055 => X"7B",  -- 123
        9056 => X"7B",  -- 123
        9057 => X"86",  -- 134
        9058 => X"7F",  -- 127
        9059 => X"84",  -- 132
        9060 => X"8B",  -- 139
        9061 => X"82",  -- 130
        9062 => X"81",  -- 129
        9063 => X"80",  -- 128
        9064 => X"79",  -- 121
        9065 => X"63",  -- 99
        9066 => X"73",  -- 115
        9067 => X"6E",  -- 110
        9068 => X"79",  -- 121
        9069 => X"70",  -- 112
        9070 => X"6C",  -- 108
        9071 => X"67",  -- 103
        9072 => X"6F",  -- 111
        9073 => X"62",  -- 98
        9074 => X"38",  -- 56
        9075 => X"30",  -- 48
        9076 => X"28",  -- 40
        9077 => X"40",  -- 64
        9078 => X"44",  -- 68
        9079 => X"3A",  -- 58
        9080 => X"57",  -- 87
        9081 => X"6C",  -- 108
        9082 => X"69",  -- 105
        9083 => X"6D",  -- 109
        9084 => X"75",  -- 117
        9085 => X"7C",  -- 124
        9086 => X"89",  -- 137
        9087 => X"8B",  -- 139
        9088 => X"85",  -- 133
        9089 => X"86",  -- 134
        9090 => X"82",  -- 130
        9091 => X"84",  -- 132
        9092 => X"88",  -- 136
        9093 => X"7F",  -- 127
        9094 => X"77",  -- 119
        9095 => X"7C",  -- 124
        9096 => X"81",  -- 129
        9097 => X"84",  -- 132
        9098 => X"85",  -- 133
        9099 => X"83",  -- 131
        9100 => X"86",  -- 134
        9101 => X"87",  -- 135
        9102 => X"83",  -- 131
        9103 => X"7E",  -- 126
        9104 => X"84",  -- 132
        9105 => X"87",  -- 135
        9106 => X"84",  -- 132
        9107 => X"7C",  -- 124
        9108 => X"79",  -- 121
        9109 => X"7D",  -- 125
        9110 => X"79",  -- 121
        9111 => X"72",  -- 114
        9112 => X"6D",  -- 109
        9113 => X"69",  -- 105
        9114 => X"5F",  -- 95
        9115 => X"56",  -- 86
        9116 => X"5A",  -- 90
        9117 => X"67",  -- 103
        9118 => X"6E",  -- 110
        9119 => X"6E",  -- 110
        9120 => X"71",  -- 113
        9121 => X"6C",  -- 108
        9122 => X"5E",  -- 94
        9123 => X"4B",  -- 75
        9124 => X"3F",  -- 63
        9125 => X"3B",  -- 59
        9126 => X"3A",  -- 58
        9127 => X"38",  -- 56
        9128 => X"3A",  -- 58
        9129 => X"3D",  -- 61
        9130 => X"45",  -- 69
        9131 => X"4A",  -- 74
        9132 => X"52",  -- 82
        9133 => X"59",  -- 89
        9134 => X"5D",  -- 93
        9135 => X"5E",  -- 94
        9136 => X"5F",  -- 95
        9137 => X"5D",  -- 93
        9138 => X"60",  -- 96
        9139 => X"6A",  -- 106
        9140 => X"6F",  -- 111
        9141 => X"6B",  -- 107
        9142 => X"65",  -- 101
        9143 => X"63",  -- 99
        9144 => X"6D",  -- 109
        9145 => X"6C",  -- 108
        9146 => X"6C",  -- 108
        9147 => X"6B",  -- 107
        9148 => X"6C",  -- 108
        9149 => X"6E",  -- 110
        9150 => X"72",  -- 114
        9151 => X"74",  -- 116
        9152 => X"6F",  -- 111
        9153 => X"72",  -- 114
        9154 => X"76",  -- 118
        9155 => X"75",  -- 117
        9156 => X"72",  -- 114
        9157 => X"71",  -- 113
        9158 => X"73",  -- 115
        9159 => X"76",  -- 118
        9160 => X"73",  -- 115
        9161 => X"78",  -- 120
        9162 => X"7E",  -- 126
        9163 => X"82",  -- 130
        9164 => X"85",  -- 133
        9165 => X"88",  -- 136
        9166 => X"8C",  -- 140
        9167 => X"8D",  -- 141
        9168 => X"8F",  -- 143
        9169 => X"8F",  -- 143
        9170 => X"95",  -- 149
        9171 => X"9F",  -- 159
        9172 => X"A2",  -- 162
        9173 => X"9F",  -- 159
        9174 => X"9F",  -- 159
        9175 => X"A4",  -- 164
        9176 => X"AC",  -- 172
        9177 => X"AD",  -- 173
        9178 => X"AF",  -- 175
        9179 => X"AF",  -- 175
        9180 => X"B0",  -- 176
        9181 => X"B1",  -- 177
        9182 => X"B4",  -- 180
        9183 => X"B6",  -- 182
        9184 => X"B6",  -- 182
        9185 => X"B1",  -- 177
        9186 => X"AE",  -- 174
        9187 => X"AC",  -- 172
        9188 => X"A6",  -- 166
        9189 => X"9D",  -- 157
        9190 => X"9E",  -- 158
        9191 => X"A6",  -- 166
        9192 => X"A1",  -- 161
        9193 => X"A1",  -- 161
        9194 => X"A5",  -- 165
        9195 => X"A6",  -- 166
        9196 => X"A2",  -- 162
        9197 => X"A2",  -- 162
        9198 => X"A5",  -- 165
        9199 => X"AA",  -- 170
        9200 => X"A6",  -- 166
        9201 => X"A4",  -- 164
        9202 => X"A4",  -- 164
        9203 => X"A5",  -- 165
        9204 => X"A5",  -- 165
        9205 => X"A3",  -- 163
        9206 => X"A0",  -- 160
        9207 => X"9D",  -- 157
        9208 => X"A2",  -- 162
        9209 => X"A1",  -- 161
        9210 => X"A2",  -- 162
        9211 => X"A6",  -- 166
        9212 => X"AB",  -- 171
        9213 => X"AD",  -- 173
        9214 => X"AB",  -- 171
        9215 => X"A8",  -- 168
        9216 => X"AA",  -- 170
        9217 => X"AB",  -- 171
        9218 => X"AC",  -- 172
        9219 => X"AC",  -- 172
        9220 => X"AF",  -- 175
        9221 => X"AF",  -- 175
        9222 => X"A9",  -- 169
        9223 => X"A0",  -- 160
        9224 => X"A0",  -- 160
        9225 => X"A1",  -- 161
        9226 => X"9E",  -- 158
        9227 => X"99",  -- 153
        9228 => X"97",  -- 151
        9229 => X"92",  -- 146
        9230 => X"7A",  -- 122
        9231 => X"61",  -- 97
        9232 => X"46",  -- 70
        9233 => X"50",  -- 80
        9234 => X"5C",  -- 92
        9235 => X"69",  -- 105
        9236 => X"7C",  -- 124
        9237 => X"92",  -- 146
        9238 => X"9E",  -- 158
        9239 => X"9E",  -- 158
        9240 => X"A7",  -- 167
        9241 => X"A6",  -- 166
        9242 => X"A6",  -- 166
        9243 => X"A6",  -- 166
        9244 => X"A5",  -- 165
        9245 => X"A3",  -- 163
        9246 => X"A1",  -- 161
        9247 => X"9D",  -- 157
        9248 => X"A6",  -- 166
        9249 => X"A6",  -- 166
        9250 => X"A2",  -- 162
        9251 => X"9C",  -- 156
        9252 => X"91",  -- 145
        9253 => X"7D",  -- 125
        9254 => X"67",  -- 103
        9255 => X"59",  -- 89
        9256 => X"5F",  -- 95
        9257 => X"61",  -- 97
        9258 => X"71",  -- 113
        9259 => X"8B",  -- 139
        9260 => X"A1",  -- 161
        9261 => X"AC",  -- 172
        9262 => X"B0",  -- 176
        9263 => X"B3",  -- 179
        9264 => X"B0",  -- 176
        9265 => X"B0",  -- 176
        9266 => X"AF",  -- 175
        9267 => X"AD",  -- 173
        9268 => X"AA",  -- 170
        9269 => X"A7",  -- 167
        9270 => X"A7",  -- 167
        9271 => X"A6",  -- 166
        9272 => X"B1",  -- 177
        9273 => X"B8",  -- 184
        9274 => X"B5",  -- 181
        9275 => X"A7",  -- 167
        9276 => X"A4",  -- 164
        9277 => X"A8",  -- 168
        9278 => X"AB",  -- 171
        9279 => X"AE",  -- 174
        9280 => X"3B",  -- 59
        9281 => X"3B",  -- 59
        9282 => X"3B",  -- 59
        9283 => X"3C",  -- 60
        9284 => X"3D",  -- 61
        9285 => X"3E",  -- 62
        9286 => X"40",  -- 64
        9287 => X"40",  -- 64
        9288 => X"40",  -- 64
        9289 => X"41",  -- 65
        9290 => X"41",  -- 65
        9291 => X"42",  -- 66
        9292 => X"42",  -- 66
        9293 => X"41",  -- 65
        9294 => X"41",  -- 65
        9295 => X"40",  -- 64
        9296 => X"40",  -- 64
        9297 => X"40",  -- 64
        9298 => X"3F",  -- 63
        9299 => X"3F",  -- 63
        9300 => X"3F",  -- 63
        9301 => X"3F",  -- 63
        9302 => X"3E",  -- 62
        9303 => X"3E",  -- 62
        9304 => X"3D",  -- 61
        9305 => X"3D",  -- 61
        9306 => X"3D",  -- 61
        9307 => X"3D",  -- 61
        9308 => X"3C",  -- 60
        9309 => X"3C",  -- 60
        9310 => X"3C",  -- 60
        9311 => X"3C",  -- 60
        9312 => X"3C",  -- 60
        9313 => X"3B",  -- 59
        9314 => X"39",  -- 57
        9315 => X"37",  -- 55
        9316 => X"37",  -- 55
        9317 => X"36",  -- 54
        9318 => X"35",  -- 53
        9319 => X"35",  -- 53
        9320 => X"32",  -- 50
        9321 => X"34",  -- 52
        9322 => X"38",  -- 56
        9323 => X"3C",  -- 60
        9324 => X"40",  -- 64
        9325 => X"47",  -- 71
        9326 => X"4F",  -- 79
        9327 => X"55",  -- 85
        9328 => X"5B",  -- 91
        9329 => X"63",  -- 99
        9330 => X"6F",  -- 111
        9331 => X"77",  -- 119
        9332 => X"79",  -- 121
        9333 => X"76",  -- 118
        9334 => X"73",  -- 115
        9335 => X"6F",  -- 111
        9336 => X"6E",  -- 110
        9337 => X"6E",  -- 110
        9338 => X"6F",  -- 111
        9339 => X"71",  -- 113
        9340 => X"74",  -- 116
        9341 => X"78",  -- 120
        9342 => X"7D",  -- 125
        9343 => X"81",  -- 129
        9344 => X"87",  -- 135
        9345 => X"85",  -- 133
        9346 => X"82",  -- 130
        9347 => X"81",  -- 129
        9348 => X"85",  -- 133
        9349 => X"88",  -- 136
        9350 => X"8C",  -- 140
        9351 => X"90",  -- 144
        9352 => X"83",  -- 131
        9353 => X"7E",  -- 126
        9354 => X"89",  -- 137
        9355 => X"8E",  -- 142
        9356 => X"7C",  -- 124
        9357 => X"70",  -- 112
        9358 => X"6A",  -- 106
        9359 => X"5B",  -- 91
        9360 => X"4B",  -- 75
        9361 => X"3B",  -- 59
        9362 => X"37",  -- 55
        9363 => X"32",  -- 50
        9364 => X"43",  -- 67
        9365 => X"41",  -- 65
        9366 => X"46",  -- 70
        9367 => X"42",  -- 66
        9368 => X"30",  -- 48
        9369 => X"33",  -- 51
        9370 => X"2D",  -- 45
        9371 => X"32",  -- 50
        9372 => X"36",  -- 54
        9373 => X"4F",  -- 79
        9374 => X"5B",  -- 91
        9375 => X"62",  -- 98
        9376 => X"6F",  -- 111
        9377 => X"82",  -- 130
        9378 => X"7A",  -- 122
        9379 => X"7B",  -- 123
        9380 => X"7C",  -- 124
        9381 => X"69",  -- 105
        9382 => X"63",  -- 99
        9383 => X"69",  -- 105
        9384 => X"67",  -- 103
        9385 => X"54",  -- 84
        9386 => X"5B",  -- 91
        9387 => X"59",  -- 89
        9388 => X"56",  -- 86
        9389 => X"50",  -- 80
        9390 => X"47",  -- 71
        9391 => X"44",  -- 68
        9392 => X"4C",  -- 76
        9393 => X"43",  -- 67
        9394 => X"2F",  -- 47
        9395 => X"2D",  -- 45
        9396 => X"2E",  -- 46
        9397 => X"38",  -- 56
        9398 => X"2E",  -- 46
        9399 => X"25",  -- 37
        9400 => X"3F",  -- 63
        9401 => X"56",  -- 86
        9402 => X"55",  -- 85
        9403 => X"5D",  -- 93
        9404 => X"6C",  -- 108
        9405 => X"79",  -- 121
        9406 => X"89",  -- 137
        9407 => X"8A",  -- 138
        9408 => X"86",  -- 134
        9409 => X"86",  -- 134
        9410 => X"87",  -- 135
        9411 => X"8B",  -- 139
        9412 => X"8C",  -- 140
        9413 => X"7E",  -- 126
        9414 => X"77",  -- 119
        9415 => X"7F",  -- 127
        9416 => X"7F",  -- 127
        9417 => X"81",  -- 129
        9418 => X"82",  -- 130
        9419 => X"81",  -- 129
        9420 => X"84",  -- 132
        9421 => X"88",  -- 136
        9422 => X"87",  -- 135
        9423 => X"83",  -- 131
        9424 => X"85",  -- 133
        9425 => X"88",  -- 136
        9426 => X"84",  -- 132
        9427 => X"7F",  -- 127
        9428 => X"80",  -- 128
        9429 => X"84",  -- 132
        9430 => X"83",  -- 131
        9431 => X"7E",  -- 126
        9432 => X"76",  -- 118
        9433 => X"73",  -- 115
        9434 => X"70",  -- 112
        9435 => X"6F",  -- 111
        9436 => X"75",  -- 117
        9437 => X"7E",  -- 126
        9438 => X"80",  -- 128
        9439 => X"7C",  -- 124
        9440 => X"6E",  -- 110
        9441 => X"5E",  -- 94
        9442 => X"47",  -- 71
        9443 => X"34",  -- 52
        9444 => X"30",  -- 48
        9445 => X"36",  -- 54
        9446 => X"35",  -- 53
        9447 => X"32",  -- 50
        9448 => X"35",  -- 53
        9449 => X"44",  -- 68
        9450 => X"53",  -- 83
        9451 => X"55",  -- 85
        9452 => X"52",  -- 82
        9453 => X"52",  -- 82
        9454 => X"59",  -- 89
        9455 => X"5D",  -- 93
        9456 => X"56",  -- 86
        9457 => X"58",  -- 88
        9458 => X"5D",  -- 93
        9459 => X"61",  -- 97
        9460 => X"60",  -- 96
        9461 => X"5E",  -- 94
        9462 => X"66",  -- 102
        9463 => X"73",  -- 115
        9464 => X"73",  -- 115
        9465 => X"71",  -- 113
        9466 => X"6F",  -- 111
        9467 => X"6D",  -- 109
        9468 => X"6C",  -- 108
        9469 => X"6C",  -- 108
        9470 => X"6D",  -- 109
        9471 => X"6E",  -- 110
        9472 => X"6A",  -- 106
        9473 => X"6D",  -- 109
        9474 => X"71",  -- 113
        9475 => X"73",  -- 115
        9476 => X"73",  -- 115
        9477 => X"73",  -- 115
        9478 => X"74",  -- 116
        9479 => X"74",  -- 116
        9480 => X"78",  -- 120
        9481 => X"7D",  -- 125
        9482 => X"81",  -- 129
        9483 => X"82",  -- 130
        9484 => X"86",  -- 134
        9485 => X"8B",  -- 139
        9486 => X"8E",  -- 142
        9487 => X"8F",  -- 143
        9488 => X"8D",  -- 141
        9489 => X"8E",  -- 142
        9490 => X"93",  -- 147
        9491 => X"9A",  -- 154
        9492 => X"9C",  -- 156
        9493 => X"9B",  -- 155
        9494 => X"9B",  -- 155
        9495 => X"9D",  -- 157
        9496 => X"AA",  -- 170
        9497 => X"AC",  -- 172
        9498 => X"AD",  -- 173
        9499 => X"AE",  -- 174
        9500 => X"AE",  -- 174
        9501 => X"B0",  -- 176
        9502 => X"B2",  -- 178
        9503 => X"B4",  -- 180
        9504 => X"B4",  -- 180
        9505 => X"B1",  -- 177
        9506 => X"B1",  -- 177
        9507 => X"AF",  -- 175
        9508 => X"AC",  -- 172
        9509 => X"A7",  -- 167
        9510 => X"A8",  -- 168
        9511 => X"AA",  -- 170
        9512 => X"A0",  -- 160
        9513 => X"9F",  -- 159
        9514 => X"A0",  -- 160
        9515 => X"A0",  -- 160
        9516 => X"A1",  -- 161
        9517 => X"A2",  -- 162
        9518 => X"A3",  -- 163
        9519 => X"A5",  -- 165
        9520 => X"A5",  -- 165
        9521 => X"A3",  -- 163
        9522 => X"A5",  -- 165
        9523 => X"A7",  -- 167
        9524 => X"A6",  -- 166
        9525 => X"A3",  -- 163
        9526 => X"A2",  -- 162
        9527 => X"A3",  -- 163
        9528 => X"A8",  -- 168
        9529 => X"A4",  -- 164
        9530 => X"A1",  -- 161
        9531 => X"A3",  -- 163
        9532 => X"A7",  -- 167
        9533 => X"A9",  -- 169
        9534 => X"A7",  -- 167
        9535 => X"A4",  -- 164
        9536 => X"9E",  -- 158
        9537 => X"A4",  -- 164
        9538 => X"AA",  -- 170
        9539 => X"AF",  -- 175
        9540 => X"B4",  -- 180
        9541 => X"B5",  -- 181
        9542 => X"AE",  -- 174
        9543 => X"A5",  -- 165
        9544 => X"A3",  -- 163
        9545 => X"A3",  -- 163
        9546 => X"9D",  -- 157
        9547 => X"96",  -- 150
        9548 => X"97",  -- 151
        9549 => X"96",  -- 150
        9550 => X"88",  -- 136
        9551 => X"76",  -- 118
        9552 => X"4C",  -- 76
        9553 => X"4A",  -- 74
        9554 => X"4B",  -- 75
        9555 => X"57",  -- 87
        9556 => X"70",  -- 112
        9557 => X"8B",  -- 139
        9558 => X"9B",  -- 155
        9559 => X"9F",  -- 159
        9560 => X"A7",  -- 167
        9561 => X"A5",  -- 165
        9562 => X"A2",  -- 162
        9563 => X"9F",  -- 159
        9564 => X"A1",  -- 161
        9565 => X"A3",  -- 163
        9566 => X"A6",  -- 166
        9567 => X"A5",  -- 165
        9568 => X"A7",  -- 167
        9569 => X"A8",  -- 168
        9570 => X"A6",  -- 166
        9571 => X"A0",  -- 160
        9572 => X"90",  -- 144
        9573 => X"7C",  -- 124
        9574 => X"68",  -- 104
        9575 => X"5C",  -- 92
        9576 => X"5A",  -- 90
        9577 => X"5D",  -- 93
        9578 => X"6E",  -- 110
        9579 => X"8B",  -- 139
        9580 => X"A2",  -- 162
        9581 => X"AE",  -- 174
        9582 => X"B5",  -- 181
        9583 => X"BA",  -- 186
        9584 => X"BA",  -- 186
        9585 => X"B6",  -- 182
        9586 => X"B0",  -- 176
        9587 => X"AC",  -- 172
        9588 => X"AA",  -- 170
        9589 => X"AD",  -- 173
        9590 => X"B1",  -- 177
        9591 => X"B3",  -- 179
        9592 => X"B7",  -- 183
        9593 => X"C0",  -- 192
        9594 => X"B4",  -- 180
        9595 => X"A4",  -- 164
        9596 => X"A7",  -- 167
        9597 => X"AE",  -- 174
        9598 => X"AF",  -- 175
        9599 => X"B1",  -- 177
        9600 => X"3B",  -- 59
        9601 => X"3B",  -- 59
        9602 => X"3B",  -- 59
        9603 => X"3C",  -- 60
        9604 => X"3D",  -- 61
        9605 => X"3E",  -- 62
        9606 => X"40",  -- 64
        9607 => X"41",  -- 65
        9608 => X"41",  -- 65
        9609 => X"41",  -- 65
        9610 => X"42",  -- 66
        9611 => X"42",  -- 66
        9612 => X"42",  -- 66
        9613 => X"42",  -- 66
        9614 => X"41",  -- 65
        9615 => X"41",  -- 65
        9616 => X"40",  -- 64
        9617 => X"40",  -- 64
        9618 => X"40",  -- 64
        9619 => X"3F",  -- 63
        9620 => X"3F",  -- 63
        9621 => X"3F",  -- 63
        9622 => X"3F",  -- 63
        9623 => X"3F",  -- 63
        9624 => X"3D",  -- 61
        9625 => X"3D",  -- 61
        9626 => X"3D",  -- 61
        9627 => X"3C",  -- 60
        9628 => X"3C",  -- 60
        9629 => X"3C",  -- 60
        9630 => X"3C",  -- 60
        9631 => X"3C",  -- 60
        9632 => X"3C",  -- 60
        9633 => X"3B",  -- 59
        9634 => X"3A",  -- 58
        9635 => X"39",  -- 57
        9636 => X"39",  -- 57
        9637 => X"39",  -- 57
        9638 => X"39",  -- 57
        9639 => X"3B",  -- 59
        9640 => X"3C",  -- 60
        9641 => X"42",  -- 66
        9642 => X"4C",  -- 76
        9643 => X"53",  -- 83
        9644 => X"58",  -- 88
        9645 => X"5E",  -- 94
        9646 => X"65",  -- 101
        9647 => X"6C",  -- 108
        9648 => X"71",  -- 113
        9649 => X"77",  -- 119
        9650 => X"81",  -- 129
        9651 => X"85",  -- 133
        9652 => X"85",  -- 133
        9653 => X"7F",  -- 127
        9654 => X"76",  -- 118
        9655 => X"71",  -- 113
        9656 => X"6B",  -- 107
        9657 => X"6C",  -- 108
        9658 => X"6B",  -- 107
        9659 => X"68",  -- 104
        9660 => X"67",  -- 103
        9661 => X"6A",  -- 106
        9662 => X"73",  -- 115
        9663 => X"79",  -- 121
        9664 => X"80",  -- 128
        9665 => X"7F",  -- 127
        9666 => X"7C",  -- 124
        9667 => X"7B",  -- 123
        9668 => X"80",  -- 128
        9669 => X"85",  -- 133
        9670 => X"89",  -- 137
        9671 => X"8A",  -- 138
        9672 => X"81",  -- 129
        9673 => X"6F",  -- 111
        9674 => X"79",  -- 121
        9675 => X"7F",  -- 127
        9676 => X"64",  -- 100
        9677 => X"55",  -- 85
        9678 => X"56",  -- 86
        9679 => X"4E",  -- 78
        9680 => X"36",  -- 54
        9681 => X"2B",  -- 43
        9682 => X"2E",  -- 46
        9683 => X"2A",  -- 42
        9684 => X"38",  -- 56
        9685 => X"33",  -- 51
        9686 => X"3C",  -- 60
        9687 => X"3D",  -- 61
        9688 => X"2F",  -- 47
        9689 => X"31",  -- 49
        9690 => X"27",  -- 39
        9691 => X"2F",  -- 47
        9692 => X"29",  -- 41
        9693 => X"3B",  -- 59
        9694 => X"3E",  -- 62
        9695 => X"47",  -- 71
        9696 => X"57",  -- 87
        9697 => X"71",  -- 113
        9698 => X"6B",  -- 107
        9699 => X"67",  -- 103
        9700 => X"61",  -- 97
        9701 => X"45",  -- 69
        9702 => X"3E",  -- 62
        9703 => X"4A",  -- 74
        9704 => X"4D",  -- 77
        9705 => X"3E",  -- 62
        9706 => X"43",  -- 67
        9707 => X"44",  -- 68
        9708 => X"34",  -- 52
        9709 => X"34",  -- 52
        9710 => X"28",  -- 40
        9711 => X"2C",  -- 44
        9712 => X"3A",  -- 58
        9713 => X"38",  -- 56
        9714 => X"3E",  -- 62
        9715 => X"3A",  -- 58
        9716 => X"3F",  -- 63
        9717 => X"31",  -- 49
        9718 => X"28",  -- 40
        9719 => X"28",  -- 40
        9720 => X"37",  -- 55
        9721 => X"49",  -- 73
        9722 => X"43",  -- 67
        9723 => X"47",  -- 71
        9724 => X"58",  -- 88
        9725 => X"67",  -- 103
        9726 => X"79",  -- 121
        9727 => X"79",  -- 121
        9728 => X"79",  -- 121
        9729 => X"83",  -- 131
        9730 => X"84",  -- 132
        9731 => X"84",  -- 132
        9732 => X"84",  -- 132
        9733 => X"7E",  -- 126
        9734 => X"7B",  -- 123
        9735 => X"83",  -- 131
        9736 => X"7B",  -- 123
        9737 => X"7F",  -- 127
        9738 => X"7F",  -- 127
        9739 => X"7E",  -- 126
        9740 => X"7F",  -- 127
        9741 => X"84",  -- 132
        9742 => X"85",  -- 133
        9743 => X"84",  -- 132
        9744 => X"88",  -- 136
        9745 => X"88",  -- 136
        9746 => X"84",  -- 132
        9747 => X"83",  -- 131
        9748 => X"83",  -- 131
        9749 => X"84",  -- 132
        9750 => X"84",  -- 132
        9751 => X"81",  -- 129
        9752 => X"81",  -- 129
        9753 => X"83",  -- 131
        9754 => X"86",  -- 134
        9755 => X"8A",  -- 138
        9756 => X"8A",  -- 138
        9757 => X"87",  -- 135
        9758 => X"88",  -- 136
        9759 => X"8B",  -- 139
        9760 => X"8A",  -- 138
        9761 => X"79",  -- 121
        9762 => X"62",  -- 98
        9763 => X"5A",  -- 90
        9764 => X"64",  -- 100
        9765 => X"6D",  -- 109
        9766 => X"6A",  -- 106
        9767 => X"60",  -- 96
        9768 => X"48",  -- 72
        9769 => X"4C",  -- 76
        9770 => X"54",  -- 84
        9771 => X"5B",  -- 91
        9772 => X"59",  -- 89
        9773 => X"54",  -- 84
        9774 => X"55",  -- 85
        9775 => X"5A",  -- 90
        9776 => X"53",  -- 83
        9777 => X"58",  -- 88
        9778 => X"5A",  -- 90
        9779 => X"57",  -- 87
        9780 => X"58",  -- 88
        9781 => X"60",  -- 96
        9782 => X"6D",  -- 109
        9783 => X"78",  -- 120
        9784 => X"70",  -- 112
        9785 => X"6F",  -- 111
        9786 => X"6D",  -- 109
        9787 => X"6C",  -- 108
        9788 => X"6C",  -- 108
        9789 => X"6B",  -- 107
        9790 => X"6B",  -- 107
        9791 => X"6A",  -- 106
        9792 => X"6F",  -- 111
        9793 => X"6E",  -- 110
        9794 => X"6E",  -- 110
        9795 => X"70",  -- 112
        9796 => X"73",  -- 115
        9797 => X"75",  -- 117
        9798 => X"76",  -- 118
        9799 => X"75",  -- 117
        9800 => X"7F",  -- 127
        9801 => X"83",  -- 131
        9802 => X"85",  -- 133
        9803 => X"83",  -- 131
        9804 => X"85",  -- 133
        9805 => X"8A",  -- 138
        9806 => X"8C",  -- 140
        9807 => X"8A",  -- 138
        9808 => X"8B",  -- 139
        9809 => X"91",  -- 145
        9810 => X"95",  -- 149
        9811 => X"94",  -- 148
        9812 => X"92",  -- 146
        9813 => X"96",  -- 150
        9814 => X"9C",  -- 156
        9815 => X"9E",  -- 158
        9816 => X"A7",  -- 167
        9817 => X"A8",  -- 168
        9818 => X"AA",  -- 170
        9819 => X"AB",  -- 171
        9820 => X"AB",  -- 171
        9821 => X"AC",  -- 172
        9822 => X"AE",  -- 174
        9823 => X"B0",  -- 176
        9824 => X"AE",  -- 174
        9825 => X"B1",  -- 177
        9826 => X"B2",  -- 178
        9827 => X"AF",  -- 175
        9828 => X"AF",  -- 175
        9829 => X"AE",  -- 174
        9830 => X"AB",  -- 171
        9831 => X"A5",  -- 165
        9832 => X"9E",  -- 158
        9833 => X"9F",  -- 159
        9834 => X"9F",  -- 159
        9835 => X"9F",  -- 159
        9836 => X"9F",  -- 159
        9837 => X"A1",  -- 161
        9838 => X"A3",  -- 163
        9839 => X"A4",  -- 164
        9840 => X"A5",  -- 165
        9841 => X"A4",  -- 164
        9842 => X"A7",  -- 167
        9843 => X"A8",  -- 168
        9844 => X"A4",  -- 164
        9845 => X"9F",  -- 159
        9846 => X"9F",  -- 159
        9847 => X"A4",  -- 164
        9848 => X"AB",  -- 171
        9849 => X"A6",  -- 166
        9850 => X"A0",  -- 160
        9851 => X"A0",  -- 160
        9852 => X"A4",  -- 164
        9853 => X"A7",  -- 167
        9854 => X"A7",  -- 167
        9855 => X"A4",  -- 164
        9856 => X"9C",  -- 156
        9857 => X"A3",  -- 163
        9858 => X"AB",  -- 171
        9859 => X"AF",  -- 175
        9860 => X"B3",  -- 179
        9861 => X"B6",  -- 182
        9862 => X"B4",  -- 180
        9863 => X"AF",  -- 175
        9864 => X"A1",  -- 161
        9865 => X"A1",  -- 161
        9866 => X"9E",  -- 158
        9867 => X"97",  -- 151
        9868 => X"92",  -- 146
        9869 => X"91",  -- 145
        9870 => X"89",  -- 137
        9871 => X"7D",  -- 125
        9872 => X"62",  -- 98
        9873 => X"50",  -- 80
        9874 => X"41",  -- 65
        9875 => X"48",  -- 72
        9876 => X"61",  -- 97
        9877 => X"7E",  -- 126
        9878 => X"92",  -- 146
        9879 => X"9C",  -- 156
        9880 => X"A0",  -- 160
        9881 => X"9E",  -- 158
        9882 => X"9B",  -- 155
        9883 => X"9B",  -- 155
        9884 => X"9D",  -- 157
        9885 => X"A1",  -- 161
        9886 => X"A4",  -- 164
        9887 => X"A4",  -- 164
        9888 => X"A2",  -- 162
        9889 => X"A2",  -- 162
        9890 => X"A3",  -- 163
        9891 => X"A1",  -- 161
        9892 => X"98",  -- 152
        9893 => X"88",  -- 136
        9894 => X"73",  -- 115
        9895 => X"67",  -- 103
        9896 => X"59",  -- 89
        9897 => X"56",  -- 86
        9898 => X"64",  -- 100
        9899 => X"82",  -- 130
        9900 => X"9F",  -- 159
        9901 => X"AE",  -- 174
        9902 => X"B4",  -- 180
        9903 => X"B9",  -- 185
        9904 => X"BB",  -- 187
        9905 => X"B7",  -- 183
        9906 => X"B3",  -- 179
        9907 => X"B0",  -- 176
        9908 => X"AF",  -- 175
        9909 => X"B2",  -- 178
        9910 => X"B5",  -- 181
        9911 => X"B6",  -- 182
        9912 => X"B7",  -- 183
        9913 => X"C3",  -- 195
        9914 => X"B7",  -- 183
        9915 => X"A7",  -- 167
        9916 => X"AE",  -- 174
        9917 => X"B3",  -- 179
        9918 => X"AD",  -- 173
        9919 => X"AD",  -- 173
        9920 => X"3B",  -- 59
        9921 => X"3A",  -- 58
        9922 => X"3C",  -- 60
        9923 => X"3C",  -- 60
        9924 => X"3D",  -- 61
        9925 => X"3F",  -- 63
        9926 => X"40",  -- 64
        9927 => X"41",  -- 65
        9928 => X"41",  -- 65
        9929 => X"41",  -- 65
        9930 => X"42",  -- 66
        9931 => X"42",  -- 66
        9932 => X"42",  -- 66
        9933 => X"42",  -- 66
        9934 => X"41",  -- 65
        9935 => X"41",  -- 65
        9936 => X"41",  -- 65
        9937 => X"41",  -- 65
        9938 => X"41",  -- 65
        9939 => X"40",  -- 64
        9940 => X"3F",  -- 63
        9941 => X"3F",  -- 63
        9942 => X"3F",  -- 63
        9943 => X"3F",  -- 63
        9944 => X"3D",  -- 61
        9945 => X"3D",  -- 61
        9946 => X"3D",  -- 61
        9947 => X"3C",  -- 60
        9948 => X"3C",  -- 60
        9949 => X"3C",  -- 60
        9950 => X"3C",  -- 60
        9951 => X"3B",  -- 59
        9952 => X"3A",  -- 58
        9953 => X"39",  -- 57
        9954 => X"39",  -- 57
        9955 => X"3A",  -- 58
        9956 => X"3E",  -- 62
        9957 => X"3F",  -- 63
        9958 => X"43",  -- 67
        9959 => X"44",  -- 68
        9960 => X"48",  -- 72
        9961 => X"52",  -- 82
        9962 => X"5F",  -- 95
        9963 => X"68",  -- 104
        9964 => X"6D",  -- 109
        9965 => X"70",  -- 112
        9966 => X"74",  -- 116
        9967 => X"78",  -- 120
        9968 => X"7B",  -- 123
        9969 => X"80",  -- 128
        9970 => X"87",  -- 135
        9971 => X"8B",  -- 139
        9972 => X"89",  -- 137
        9973 => X"83",  -- 131
        9974 => X"7D",  -- 125
        9975 => X"78",  -- 120
        9976 => X"76",  -- 118
        9977 => X"73",  -- 115
        9978 => X"6D",  -- 109
        9979 => X"63",  -- 99
        9980 => X"5E",  -- 94
        9981 => X"62",  -- 98
        9982 => X"6E",  -- 110
        9983 => X"78",  -- 120
        9984 => X"7A",  -- 122
        9985 => X"78",  -- 120
        9986 => X"77",  -- 119
        9987 => X"77",  -- 119
        9988 => X"79",  -- 121
        9989 => X"7D",  -- 125
        9990 => X"80",  -- 128
        9991 => X"81",  -- 129
        9992 => X"83",  -- 131
        9993 => X"67",  -- 103
        9994 => X"69",  -- 105
        9995 => X"6C",  -- 108
        9996 => X"50",  -- 80
        9997 => X"43",  -- 67
        9998 => X"4E",  -- 78
        9999 => X"51",  -- 81
        10000 => X"33",  -- 51
        10001 => X"2D",  -- 45
        10002 => X"32",  -- 50
        10003 => X"2D",  -- 45
        10004 => X"35",  -- 53
        10005 => X"2B",  -- 43
        10006 => X"35",  -- 53
        10007 => X"37",  -- 55
        10008 => X"32",  -- 50
        10009 => X"33",  -- 51
        10010 => X"29",  -- 41
        10011 => X"30",  -- 48
        10012 => X"22",  -- 34
        10013 => X"2D",  -- 45
        10014 => X"2A",  -- 42
        10015 => X"35",  -- 53
        10016 => X"38",  -- 56
        10017 => X"57",  -- 87
        10018 => X"55",  -- 85
        10019 => X"52",  -- 82
        10020 => X"4C",  -- 76
        10021 => X"2F",  -- 47
        10022 => X"2A",  -- 42
        10023 => X"3A",  -- 58
        10024 => X"32",  -- 50
        10025 => X"2B",  -- 43
        10026 => X"30",  -- 48
        10027 => X"39",  -- 57
        10028 => X"26",  -- 38
        10029 => X"2E",  -- 46
        10030 => X"25",  -- 37
        10031 => X"32",  -- 50
        10032 => X"3A",  -- 58
        10033 => X"3E",  -- 62
        10034 => X"50",  -- 80
        10035 => X"47",  -- 71
        10036 => X"48",  -- 72
        10037 => X"2E",  -- 46
        10038 => X"2A",  -- 42
        10039 => X"37",  -- 55
        10040 => X"4A",  -- 74
        10041 => X"54",  -- 84
        10042 => X"41",  -- 65
        10043 => X"38",  -- 56
        10044 => X"43",  -- 67
        10045 => X"54",  -- 84
        10046 => X"64",  -- 100
        10047 => X"65",  -- 101
        10048 => X"6B",  -- 107
        10049 => X"7C",  -- 124
        10050 => X"7F",  -- 127
        10051 => X"78",  -- 120
        10052 => X"79",  -- 121
        10053 => X"7E",  -- 126
        10054 => X"80",  -- 128
        10055 => X"83",  -- 131
        10056 => X"7F",  -- 127
        10057 => X"83",  -- 131
        10058 => X"82",  -- 130
        10059 => X"7F",  -- 127
        10060 => X"7E",  -- 126
        10061 => X"81",  -- 129
        10062 => X"84",  -- 132
        10063 => X"85",  -- 133
        10064 => X"86",  -- 134
        10065 => X"84",  -- 132
        10066 => X"83",  -- 131
        10067 => X"87",  -- 135
        10068 => X"88",  -- 136
        10069 => X"88",  -- 136
        10070 => X"87",  -- 135
        10071 => X"89",  -- 137
        10072 => X"8A",  -- 138
        10073 => X"8E",  -- 142
        10074 => X"95",  -- 149
        10075 => X"97",  -- 151
        10076 => X"8E",  -- 142
        10077 => X"85",  -- 133
        10078 => X"89",  -- 137
        10079 => X"94",  -- 148
        10080 => X"93",  -- 147
        10081 => X"93",  -- 147
        10082 => X"91",  -- 145
        10083 => X"8A",  -- 138
        10084 => X"86",  -- 134
        10085 => X"86",  -- 134
        10086 => X"88",  -- 136
        10087 => X"86",  -- 134
        10088 => X"6F",  -- 111
        10089 => X"57",  -- 87
        10090 => X"4E",  -- 78
        10091 => X"59",  -- 89
        10092 => X"60",  -- 96
        10093 => X"55",  -- 85
        10094 => X"4D",  -- 77
        10095 => X"50",  -- 80
        10096 => X"54",  -- 84
        10097 => X"59",  -- 89
        10098 => X"56",  -- 86
        10099 => X"51",  -- 81
        10100 => X"5A",  -- 90
        10101 => X"6F",  -- 111
        10102 => X"76",  -- 118
        10103 => X"71",  -- 113
        10104 => X"6D",  -- 109
        10105 => X"6D",  -- 109
        10106 => X"6C",  -- 108
        10107 => X"6D",  -- 109
        10108 => X"6F",  -- 111
        10109 => X"70",  -- 112
        10110 => X"70",  -- 112
        10111 => X"6F",  -- 111
        10112 => X"78",  -- 120
        10113 => X"74",  -- 116
        10114 => X"6F",  -- 111
        10115 => X"70",  -- 112
        10116 => X"74",  -- 116
        10117 => X"76",  -- 118
        10118 => X"77",  -- 119
        10119 => X"75",  -- 117
        10120 => X"77",  -- 119
        10121 => X"7B",  -- 123
        10122 => X"7D",  -- 125
        10123 => X"7D",  -- 125
        10124 => X"80",  -- 128
        10125 => X"87",  -- 135
        10126 => X"8A",  -- 138
        10127 => X"89",  -- 137
        10128 => X"89",  -- 137
        10129 => X"95",  -- 149
        10130 => X"98",  -- 152
        10131 => X"90",  -- 144
        10132 => X"8B",  -- 139
        10133 => X"92",  -- 146
        10134 => X"9C",  -- 156
        10135 => X"A2",  -- 162
        10136 => X"A4",  -- 164
        10137 => X"A5",  -- 165
        10138 => X"A7",  -- 167
        10139 => X"A8",  -- 168
        10140 => X"A8",  -- 168
        10141 => X"A9",  -- 169
        10142 => X"AA",  -- 170
        10143 => X"AB",  -- 171
        10144 => X"A8",  -- 168
        10145 => X"AD",  -- 173
        10146 => X"AF",  -- 175
        10147 => X"AE",  -- 174
        10148 => X"AE",  -- 174
        10149 => X"B0",  -- 176
        10150 => X"A8",  -- 168
        10151 => X"9C",  -- 156
        10152 => X"9D",  -- 157
        10153 => X"A0",  -- 160
        10154 => X"A2",  -- 162
        10155 => X"A0",  -- 160
        10156 => X"9E",  -- 158
        10157 => X"A0",  -- 160
        10158 => X"A4",  -- 164
        10159 => X"A7",  -- 167
        10160 => X"A5",  -- 165
        10161 => X"A5",  -- 165
        10162 => X"A8",  -- 168
        10163 => X"A8",  -- 168
        10164 => X"A2",  -- 162
        10165 => X"9B",  -- 155
        10166 => X"9B",  -- 155
        10167 => X"A2",  -- 162
        10168 => X"AA",  -- 170
        10169 => X"A4",  -- 164
        10170 => X"9E",  -- 158
        10171 => X"9E",  -- 158
        10172 => X"A4",  -- 164
        10173 => X"A8",  -- 168
        10174 => X"A9",  -- 169
        10175 => X"A8",  -- 168
        10176 => X"A5",  -- 165
        10177 => X"AA",  -- 170
        10178 => X"AD",  -- 173
        10179 => X"AB",  -- 171
        10180 => X"AB",  -- 171
        10181 => X"AC",  -- 172
        10182 => X"AB",  -- 171
        10183 => X"A7",  -- 167
        10184 => X"99",  -- 153
        10185 => X"9D",  -- 157
        10186 => X"9D",  -- 157
        10187 => X"9B",  -- 155
        10188 => X"97",  -- 151
        10189 => X"94",  -- 148
        10190 => X"8F",  -- 143
        10191 => X"8A",  -- 138
        10192 => X"7A",  -- 122
        10193 => X"5B",  -- 91
        10194 => X"40",  -- 64
        10195 => X"42",  -- 66
        10196 => X"57",  -- 87
        10197 => X"71",  -- 113
        10198 => X"87",  -- 135
        10199 => X"94",  -- 148
        10200 => X"9C",  -- 156
        10201 => X"9C",  -- 156
        10202 => X"9E",  -- 158
        10203 => X"A1",  -- 161
        10204 => X"A2",  -- 162
        10205 => X"A2",  -- 162
        10206 => X"A2",  -- 162
        10207 => X"9F",  -- 159
        10208 => X"9C",  -- 156
        10209 => X"9D",  -- 157
        10210 => X"9F",  -- 159
        10211 => X"A4",  -- 164
        10212 => X"A1",  -- 161
        10213 => X"95",  -- 149
        10214 => X"82",  -- 130
        10215 => X"71",  -- 113
        10216 => X"65",  -- 101
        10217 => X"5C",  -- 92
        10218 => X"61",  -- 97
        10219 => X"7D",  -- 125
        10220 => X"98",  -- 152
        10221 => X"A5",  -- 165
        10222 => X"A7",  -- 167
        10223 => X"A9",  -- 169
        10224 => X"B0",  -- 176
        10225 => X"B1",  -- 177
        10226 => X"B1",  -- 177
        10227 => X"B1",  -- 177
        10228 => X"B1",  -- 177
        10229 => X"AF",  -- 175
        10230 => X"AC",  -- 172
        10231 => X"AB",  -- 171
        10232 => X"B2",  -- 178
        10233 => X"C2",  -- 194
        10234 => X"BA",  -- 186
        10235 => X"AD",  -- 173
        10236 => X"B6",  -- 182
        10237 => X"B7",  -- 183
        10238 => X"AA",  -- 170
        10239 => X"A6",  -- 166
        10240 => X"39",  -- 57
        10241 => X"3A",  -- 58
        10242 => X"3B",  -- 59
        10243 => X"3C",  -- 60
        10244 => X"3F",  -- 63
        10245 => X"40",  -- 64
        10246 => X"42",  -- 66
        10247 => X"42",  -- 66
        10248 => X"40",  -- 64
        10249 => X"41",  -- 65
        10250 => X"41",  -- 65
        10251 => X"42",  -- 66
        10252 => X"42",  -- 66
        10253 => X"42",  -- 66
        10254 => X"40",  -- 64
        10255 => X"41",  -- 65
        10256 => X"44",  -- 68
        10257 => X"42",  -- 66
        10258 => X"40",  -- 64
        10259 => X"3D",  -- 61
        10260 => X"3C",  -- 60
        10261 => X"3D",  -- 61
        10262 => X"3E",  -- 62
        10263 => X"3F",  -- 63
        10264 => X"3C",  -- 60
        10265 => X"3C",  -- 60
        10266 => X"3C",  -- 60
        10267 => X"3D",  -- 61
        10268 => X"3D",  -- 61
        10269 => X"3C",  -- 60
        10270 => X"3B",  -- 59
        10271 => X"3A",  -- 58
        10272 => X"39",  -- 57
        10273 => X"3B",  -- 59
        10274 => X"3C",  -- 60
        10275 => X"41",  -- 65
        10276 => X"4B",  -- 75
        10277 => X"58",  -- 88
        10278 => X"5B",  -- 91
        10279 => X"58",  -- 88
        10280 => X"61",  -- 97
        10281 => X"6B",  -- 107
        10282 => X"74",  -- 116
        10283 => X"79",  -- 121
        10284 => X"79",  -- 121
        10285 => X"79",  -- 121
        10286 => X"7B",  -- 123
        10287 => X"7D",  -- 125
        10288 => X"82",  -- 130
        10289 => X"85",  -- 133
        10290 => X"88",  -- 136
        10291 => X"87",  -- 135
        10292 => X"83",  -- 131
        10293 => X"80",  -- 128
        10294 => X"80",  -- 128
        10295 => X"7F",  -- 127
        10296 => X"7C",  -- 124
        10297 => X"7B",  -- 123
        10298 => X"72",  -- 114
        10299 => X"61",  -- 97
        10300 => X"59",  -- 89
        10301 => X"62",  -- 98
        10302 => X"74",  -- 116
        10303 => X"7E",  -- 126
        10304 => X"82",  -- 130
        10305 => X"7B",  -- 123
        10306 => X"78",  -- 120
        10307 => X"79",  -- 121
        10308 => X"79",  -- 121
        10309 => X"74",  -- 116
        10310 => X"74",  -- 116
        10311 => X"76",  -- 118
        10312 => X"68",  -- 104
        10313 => X"6B",  -- 107
        10314 => X"5D",  -- 93
        10315 => X"69",  -- 105
        10316 => X"49",  -- 73
        10317 => X"5B",  -- 91
        10318 => X"58",  -- 88
        10319 => X"63",  -- 99
        10320 => X"4E",  -- 78
        10321 => X"41",  -- 65
        10322 => X"40",  -- 64
        10323 => X"34",  -- 52
        10324 => X"37",  -- 55
        10325 => X"39",  -- 57
        10326 => X"2C",  -- 44
        10327 => X"3B",  -- 59
        10328 => X"2B",  -- 43
        10329 => X"2E",  -- 46
        10330 => X"2A",  -- 42
        10331 => X"26",  -- 38
        10332 => X"27",  -- 39
        10333 => X"20",  -- 32
        10334 => X"1C",  -- 28
        10335 => X"23",  -- 35
        10336 => X"38",  -- 56
        10337 => X"46",  -- 70
        10338 => X"3E",  -- 62
        10339 => X"35",  -- 53
        10340 => X"2C",  -- 44
        10341 => X"2D",  -- 45
        10342 => X"35",  -- 53
        10343 => X"2B",  -- 43
        10344 => X"28",  -- 40
        10345 => X"29",  -- 41
        10346 => X"29",  -- 41
        10347 => X"26",  -- 38
        10348 => X"22",  -- 34
        10349 => X"22",  -- 34
        10350 => X"28",  -- 40
        10351 => X"30",  -- 48
        10352 => X"32",  -- 50
        10353 => X"3D",  -- 61
        10354 => X"47",  -- 71
        10355 => X"40",  -- 64
        10356 => X"51",  -- 81
        10357 => X"52",  -- 82
        10358 => X"3F",  -- 63
        10359 => X"54",  -- 84
        10360 => X"52",  -- 82
        10361 => X"56",  -- 86
        10362 => X"5B",  -- 91
        10363 => X"59",  -- 89
        10364 => X"3A",  -- 58
        10365 => X"44",  -- 68
        10366 => X"3F",  -- 63
        10367 => X"4C",  -- 76
        10368 => X"6C",  -- 108
        10369 => X"57",  -- 87
        10370 => X"6D",  -- 109
        10371 => X"6F",  -- 111
        10372 => X"5B",  -- 91
        10373 => X"6F",  -- 111
        10374 => X"82",  -- 130
        10375 => X"7C",  -- 124
        10376 => X"77",  -- 119
        10377 => X"79",  -- 121
        10378 => X"7C",  -- 124
        10379 => X"7F",  -- 127
        10380 => X"82",  -- 130
        10381 => X"83",  -- 131
        10382 => X"83",  -- 131
        10383 => X"82",  -- 130
        10384 => X"8B",  -- 139
        10385 => X"89",  -- 137
        10386 => X"85",  -- 133
        10387 => X"85",  -- 133
        10388 => X"87",  -- 135
        10389 => X"88",  -- 136
        10390 => X"8C",  -- 140
        10391 => X"8E",  -- 142
        10392 => X"94",  -- 148
        10393 => X"97",  -- 151
        10394 => X"97",  -- 151
        10395 => X"93",  -- 147
        10396 => X"8F",  -- 143
        10397 => X"8F",  -- 143
        10398 => X"93",  -- 147
        10399 => X"9B",  -- 155
        10400 => X"9C",  -- 156
        10401 => X"9B",  -- 155
        10402 => X"9B",  -- 155
        10403 => X"9D",  -- 157
        10404 => X"A0",  -- 160
        10405 => X"9E",  -- 158
        10406 => X"9B",  -- 155
        10407 => X"95",  -- 149
        10408 => X"7C",  -- 124
        10409 => X"6E",  -- 110
        10410 => X"61",  -- 97
        10411 => X"5A",  -- 90
        10412 => X"51",  -- 81
        10413 => X"4B",  -- 75
        10414 => X"4B",  -- 75
        10415 => X"52",  -- 82
        10416 => X"55",  -- 85
        10417 => X"59",  -- 89
        10418 => X"5E",  -- 94
        10419 => X"63",  -- 99
        10420 => X"67",  -- 103
        10421 => X"69",  -- 105
        10422 => X"6E",  -- 110
        10423 => X"70",  -- 112
        10424 => X"6C",  -- 108
        10425 => X"6D",  -- 109
        10426 => X"6F",  -- 111
        10427 => X"6F",  -- 111
        10428 => X"6E",  -- 110
        10429 => X"6D",  -- 109
        10430 => X"6E",  -- 110
        10431 => X"6E",  -- 110
        10432 => X"6A",  -- 106
        10433 => X"6A",  -- 106
        10434 => X"6E",  -- 110
        10435 => X"73",  -- 115
        10436 => X"74",  -- 116
        10437 => X"75",  -- 117
        10438 => X"79",  -- 121
        10439 => X"7E",  -- 126
        10440 => X"81",  -- 129
        10441 => X"7A",  -- 122
        10442 => X"76",  -- 118
        10443 => X"7C",  -- 124
        10444 => X"84",  -- 132
        10445 => X"89",  -- 137
        10446 => X"8B",  -- 139
        10447 => X"8D",  -- 141
        10448 => X"92",  -- 146
        10449 => X"94",  -- 148
        10450 => X"95",  -- 149
        10451 => X"93",  -- 147
        10452 => X"91",  -- 145
        10453 => X"93",  -- 147
        10454 => X"99",  -- 153
        10455 => X"9E",  -- 158
        10456 => X"A4",  -- 164
        10457 => X"A8",  -- 168
        10458 => X"B1",  -- 177
        10459 => X"B7",  -- 183
        10460 => X"B0",  -- 176
        10461 => X"A5",  -- 165
        10462 => X"A8",  -- 168
        10463 => X"B3",  -- 179
        10464 => X"AE",  -- 174
        10465 => X"AF",  -- 175
        10466 => X"AE",  -- 174
        10467 => X"A9",  -- 169
        10468 => X"A6",  -- 166
        10469 => X"A3",  -- 163
        10470 => X"9D",  -- 157
        10471 => X"95",  -- 149
        10472 => X"97",  -- 151
        10473 => X"9C",  -- 156
        10474 => X"A0",  -- 160
        10475 => X"A0",  -- 160
        10476 => X"9C",  -- 156
        10477 => X"9B",  -- 155
        10478 => X"9C",  -- 156
        10479 => X"9F",  -- 159
        10480 => X"A4",  -- 164
        10481 => X"A4",  -- 164
        10482 => X"A3",  -- 163
        10483 => X"A1",  -- 161
        10484 => X"9C",  -- 156
        10485 => X"9A",  -- 154
        10486 => X"9D",  -- 157
        10487 => X"A1",  -- 161
        10488 => X"A1",  -- 161
        10489 => X"A2",  -- 162
        10490 => X"A3",  -- 163
        10491 => X"A3",  -- 163
        10492 => X"A5",  -- 165
        10493 => X"A6",  -- 166
        10494 => X"A7",  -- 167
        10495 => X"A8",  -- 168
        10496 => X"AC",  -- 172
        10497 => X"AE",  -- 174
        10498 => X"B0",  -- 176
        10499 => X"AC",  -- 172
        10500 => X"A6",  -- 166
        10501 => X"A1",  -- 161
        10502 => X"9F",  -- 159
        10503 => X"9F",  -- 159
        10504 => X"9F",  -- 159
        10505 => X"9B",  -- 155
        10506 => X"96",  -- 150
        10507 => X"95",  -- 149
        10508 => X"9A",  -- 154
        10509 => X"9B",  -- 155
        10510 => X"9B",  -- 155
        10511 => X"99",  -- 153
        10512 => X"8B",  -- 139
        10513 => X"65",  -- 101
        10514 => X"4F",  -- 79
        10515 => X"50",  -- 80
        10516 => X"52",  -- 82
        10517 => X"5E",  -- 94
        10518 => X"7A",  -- 122
        10519 => X"8F",  -- 143
        10520 => X"9A",  -- 154
        10521 => X"9D",  -- 157
        10522 => X"A0",  -- 160
        10523 => X"A1",  -- 161
        10524 => X"9F",  -- 159
        10525 => X"9E",  -- 158
        10526 => X"A3",  -- 163
        10527 => X"A8",  -- 168
        10528 => X"A0",  -- 160
        10529 => X"A4",  -- 164
        10530 => X"A7",  -- 167
        10531 => X"A8",  -- 168
        10532 => X"A3",  -- 163
        10533 => X"96",  -- 150
        10534 => X"84",  -- 132
        10535 => X"73",  -- 115
        10536 => X"5C",  -- 92
        10537 => X"5E",  -- 94
        10538 => X"67",  -- 103
        10539 => X"76",  -- 118
        10540 => X"8A",  -- 138
        10541 => X"9A",  -- 154
        10542 => X"A1",  -- 161
        10543 => X"A5",  -- 165
        10544 => X"AE",  -- 174
        10545 => X"AE",  -- 174
        10546 => X"B0",  -- 176
        10547 => X"B2",  -- 178
        10548 => X"B2",  -- 178
        10549 => X"B4",  -- 180
        10550 => X"B5",  -- 181
        10551 => X"B5",  -- 181
        10552 => X"B9",  -- 185
        10553 => X"C4",  -- 196
        10554 => X"B9",  -- 185
        10555 => X"AD",  -- 173
        10556 => X"B5",  -- 181
        10557 => X"B6",  -- 182
        10558 => X"AD",  -- 173
        10559 => X"B1",  -- 177
        10560 => X"39",  -- 57
        10561 => X"3A",  -- 58
        10562 => X"3B",  -- 59
        10563 => X"3C",  -- 60
        10564 => X"3E",  -- 62
        10565 => X"3F",  -- 63
        10566 => X"41",  -- 65
        10567 => X"42",  -- 66
        10568 => X"45",  -- 69
        10569 => X"45",  -- 69
        10570 => X"44",  -- 68
        10571 => X"44",  -- 68
        10572 => X"44",  -- 68
        10573 => X"42",  -- 66
        10574 => X"41",  -- 65
        10575 => X"41",  -- 65
        10576 => X"3E",  -- 62
        10577 => X"3D",  -- 61
        10578 => X"3D",  -- 61
        10579 => X"3E",  -- 62
        10580 => X"3E",  -- 62
        10581 => X"3D",  -- 61
        10582 => X"3D",  -- 61
        10583 => X"3F",  -- 63
        10584 => X"3F",  -- 63
        10585 => X"3D",  -- 61
        10586 => X"3C",  -- 60
        10587 => X"3C",  -- 60
        10588 => X"3E",  -- 62
        10589 => X"3F",  -- 63
        10590 => X"3F",  -- 63
        10591 => X"3F",  -- 63
        10592 => X"42",  -- 66
        10593 => X"46",  -- 70
        10594 => X"4B",  -- 75
        10595 => X"4F",  -- 79
        10596 => X"59",  -- 89
        10597 => X"64",  -- 100
        10598 => X"68",  -- 104
        10599 => X"67",  -- 103
        10600 => X"75",  -- 117
        10601 => X"79",  -- 121
        10602 => X"80",  -- 128
        10603 => X"80",  -- 128
        10604 => X"7C",  -- 124
        10605 => X"7A",  -- 122
        10606 => X"7E",  -- 126
        10607 => X"82",  -- 130
        10608 => X"87",  -- 135
        10609 => X"88",  -- 136
        10610 => X"87",  -- 135
        10611 => X"83",  -- 131
        10612 => X"7F",  -- 127
        10613 => X"7D",  -- 125
        10614 => X"80",  -- 128
        10615 => X"82",  -- 130
        10616 => X"86",  -- 134
        10617 => X"86",  -- 134
        10618 => X"7D",  -- 125
        10619 => X"70",  -- 112
        10620 => X"68",  -- 104
        10621 => X"6D",  -- 109
        10622 => X"78",  -- 120
        10623 => X"80",  -- 128
        10624 => X"7D",  -- 125
        10625 => X"79",  -- 121
        10626 => X"78",  -- 120
        10627 => X"7B",  -- 123
        10628 => X"77",  -- 119
        10629 => X"6F",  -- 111
        10630 => X"67",  -- 103
        10631 => X"67",  -- 103
        10632 => X"5C",  -- 92
        10633 => X"66",  -- 102
        10634 => X"62",  -- 98
        10635 => X"73",  -- 115
        10636 => X"5E",  -- 94
        10637 => X"6D",  -- 109
        10638 => X"5C",  -- 92
        10639 => X"54",  -- 84
        10640 => X"51",  -- 81
        10641 => X"49",  -- 73
        10642 => X"49",  -- 73
        10643 => X"42",  -- 66
        10644 => X"49",  -- 73
        10645 => X"4B",  -- 75
        10646 => X"3A",  -- 58
        10647 => X"46",  -- 70
        10648 => X"2C",  -- 44
        10649 => X"30",  -- 48
        10650 => X"26",  -- 38
        10651 => X"26",  -- 38
        10652 => X"22",  -- 34
        10653 => X"24",  -- 36
        10654 => X"1E",  -- 30
        10655 => X"25",  -- 37
        10656 => X"23",  -- 35
        10657 => X"30",  -- 48
        10658 => X"2A",  -- 42
        10659 => X"27",  -- 39
        10660 => X"25",  -- 37
        10661 => X"24",  -- 36
        10662 => X"2F",  -- 47
        10663 => X"28",  -- 40
        10664 => X"21",  -- 33
        10665 => X"1D",  -- 29
        10666 => X"1A",  -- 26
        10667 => X"1F",  -- 31
        10668 => X"25",  -- 37
        10669 => X"29",  -- 41
        10670 => X"28",  -- 40
        10671 => X"25",  -- 37
        10672 => X"2D",  -- 45
        10673 => X"30",  -- 48
        10674 => X"35",  -- 53
        10675 => X"34",  -- 52
        10676 => X"4A",  -- 74
        10677 => X"4F",  -- 79
        10678 => X"3E",  -- 62
        10679 => X"54",  -- 84
        10680 => X"63",  -- 99
        10681 => X"58",  -- 88
        10682 => X"5F",  -- 95
        10683 => X"69",  -- 105
        10684 => X"4E",  -- 78
        10685 => X"45",  -- 69
        10686 => X"38",  -- 56
        10687 => X"48",  -- 72
        10688 => X"46",  -- 70
        10689 => X"4D",  -- 77
        10690 => X"50",  -- 80
        10691 => X"3E",  -- 62
        10692 => X"4A",  -- 74
        10693 => X"6F",  -- 111
        10694 => X"78",  -- 120
        10695 => X"72",  -- 114
        10696 => X"75",  -- 117
        10697 => X"74",  -- 116
        10698 => X"7F",  -- 127
        10699 => X"8B",  -- 139
        10700 => X"8B",  -- 139
        10701 => X"80",  -- 128
        10702 => X"7A",  -- 122
        10703 => X"7E",  -- 126
        10704 => X"88",  -- 136
        10705 => X"84",  -- 132
        10706 => X"82",  -- 130
        10707 => X"82",  -- 130
        10708 => X"84",  -- 132
        10709 => X"88",  -- 136
        10710 => X"8C",  -- 140
        10711 => X"8F",  -- 143
        10712 => X"8F",  -- 143
        10713 => X"88",  -- 136
        10714 => X"85",  -- 133
        10715 => X"88",  -- 136
        10716 => X"90",  -- 144
        10717 => X"98",  -- 152
        10718 => X"9C",  -- 156
        10719 => X"9A",  -- 154
        10720 => X"A4",  -- 164
        10721 => X"A0",  -- 160
        10722 => X"9F",  -- 159
        10723 => X"A1",  -- 161
        10724 => X"A4",  -- 164
        10725 => X"A8",  -- 168
        10726 => X"A8",  -- 168
        10727 => X"A6",  -- 166
        10728 => X"97",  -- 151
        10729 => X"7F",  -- 127
        10730 => X"60",  -- 96
        10731 => X"50",  -- 80
        10732 => X"4E",  -- 78
        10733 => X"55",  -- 85
        10734 => X"60",  -- 96
        10735 => X"67",  -- 103
        10736 => X"63",  -- 99
        10737 => X"63",  -- 99
        10738 => X"63",  -- 99
        10739 => X"64",  -- 100
        10740 => X"66",  -- 102
        10741 => X"68",  -- 104
        10742 => X"6A",  -- 106
        10743 => X"6B",  -- 107
        10744 => X"70",  -- 112
        10745 => X"6C",  -- 108
        10746 => X"67",  -- 103
        10747 => X"64",  -- 100
        10748 => X"65",  -- 101
        10749 => X"69",  -- 105
        10750 => X"6F",  -- 111
        10751 => X"72",  -- 114
        10752 => X"6E",  -- 110
        10753 => X"73",  -- 115
        10754 => X"76",  -- 118
        10755 => X"75",  -- 117
        10756 => X"72",  -- 114
        10757 => X"74",  -- 116
        10758 => X"7A",  -- 122
        10759 => X"7F",  -- 127
        10760 => X"7C",  -- 124
        10761 => X"79",  -- 121
        10762 => X"78",  -- 120
        10763 => X"7B",  -- 123
        10764 => X"7F",  -- 127
        10765 => X"82",  -- 130
        10766 => X"88",  -- 136
        10767 => X"8E",  -- 142
        10768 => X"8E",  -- 142
        10769 => X"90",  -- 144
        10770 => X"91",  -- 145
        10771 => X"90",  -- 144
        10772 => X"8E",  -- 142
        10773 => X"8F",  -- 143
        10774 => X"95",  -- 149
        10775 => X"9A",  -- 154
        10776 => X"A3",  -- 163
        10777 => X"A9",  -- 169
        10778 => X"AD",  -- 173
        10779 => X"AD",  -- 173
        10780 => X"AC",  -- 172
        10781 => X"AB",  -- 171
        10782 => X"AA",  -- 170
        10783 => X"A9",  -- 169
        10784 => X"AC",  -- 172
        10785 => X"AD",  -- 173
        10786 => X"AC",  -- 172
        10787 => X"A7",  -- 167
        10788 => X"A4",  -- 164
        10789 => X"A2",  -- 162
        10790 => X"9D",  -- 157
        10791 => X"98",  -- 152
        10792 => X"9B",  -- 155
        10793 => X"9E",  -- 158
        10794 => X"A1",  -- 161
        10795 => X"A0",  -- 160
        10796 => X"9E",  -- 158
        10797 => X"9D",  -- 157
        10798 => X"9E",  -- 158
        10799 => X"A2",  -- 162
        10800 => X"A3",  -- 163
        10801 => X"A5",  -- 165
        10802 => X"A4",  -- 164
        10803 => X"9F",  -- 159
        10804 => X"9F",  -- 159
        10805 => X"A1",  -- 161
        10806 => X"A1",  -- 161
        10807 => X"9B",  -- 155
        10808 => X"98",  -- 152
        10809 => X"9C",  -- 156
        10810 => X"A0",  -- 160
        10811 => X"A4",  -- 164
        10812 => X"A8",  -- 168
        10813 => X"AB",  -- 171
        10814 => X"AE",  -- 174
        10815 => X"AD",  -- 173
        10816 => X"AA",  -- 170
        10817 => X"AC",  -- 172
        10818 => X"B0",  -- 176
        10819 => X"B0",  -- 176
        10820 => X"AB",  -- 171
        10821 => X"A6",  -- 166
        10822 => X"A2",  -- 162
        10823 => X"A1",  -- 161
        10824 => X"A2",  -- 162
        10825 => X"9D",  -- 157
        10826 => X"99",  -- 153
        10827 => X"9A",  -- 154
        10828 => X"9D",  -- 157
        10829 => X"A1",  -- 161
        10830 => X"A1",  -- 161
        10831 => X"A0",  -- 160
        10832 => X"8F",  -- 143
        10833 => X"77",  -- 119
        10834 => X"63",  -- 99
        10835 => X"55",  -- 85
        10836 => X"4C",  -- 76
        10837 => X"58",  -- 88
        10838 => X"73",  -- 115
        10839 => X"86",  -- 134
        10840 => X"96",  -- 150
        10841 => X"9C",  -- 156
        10842 => X"A2",  -- 162
        10843 => X"A3",  -- 163
        10844 => X"9F",  -- 159
        10845 => X"9C",  -- 156
        10846 => X"9F",  -- 159
        10847 => X"A2",  -- 162
        10848 => X"A3",  -- 163
        10849 => X"A3",  -- 163
        10850 => X"A1",  -- 161
        10851 => X"9D",  -- 157
        10852 => X"98",  -- 152
        10853 => X"8F",  -- 143
        10854 => X"7F",  -- 127
        10855 => X"72",  -- 114
        10856 => X"62",  -- 98
        10857 => X"65",  -- 101
        10858 => X"6D",  -- 109
        10859 => X"7A",  -- 122
        10860 => X"8B",  -- 139
        10861 => X"99",  -- 153
        10862 => X"A6",  -- 166
        10863 => X"AC",  -- 172
        10864 => X"AE",  -- 174
        10865 => X"AF",  -- 175
        10866 => X"B1",  -- 177
        10867 => X"B2",  -- 178
        10868 => X"B5",  -- 181
        10869 => X"B5",  -- 181
        10870 => X"B6",  -- 182
        10871 => X"B6",  -- 182
        10872 => X"B7",  -- 183
        10873 => X"C1",  -- 193
        10874 => X"B8",  -- 184
        10875 => X"AD",  -- 173
        10876 => X"B3",  -- 179
        10877 => X"B3",  -- 179
        10878 => X"AE",  -- 174
        10879 => X"B0",  -- 176
        10880 => X"3A",  -- 58
        10881 => X"3B",  -- 59
        10882 => X"3C",  -- 60
        10883 => X"3D",  -- 61
        10884 => X"3E",  -- 62
        10885 => X"40",  -- 64
        10886 => X"41",  -- 65
        10887 => X"41",  -- 65
        10888 => X"42",  -- 66
        10889 => X"42",  -- 66
        10890 => X"42",  -- 66
        10891 => X"42",  -- 66
        10892 => X"41",  -- 65
        10893 => X"40",  -- 64
        10894 => X"3F",  -- 63
        10895 => X"3F",  -- 63
        10896 => X"3D",  -- 61
        10897 => X"3E",  -- 62
        10898 => X"3E",  -- 62
        10899 => X"3F",  -- 63
        10900 => X"3E",  -- 62
        10901 => X"3E",  -- 62
        10902 => X"3C",  -- 60
        10903 => X"3C",  -- 60
        10904 => X"3E",  -- 62
        10905 => X"3E",  -- 62
        10906 => X"3D",  -- 61
        10907 => X"3E",  -- 62
        10908 => X"40",  -- 64
        10909 => X"44",  -- 68
        10910 => X"46",  -- 70
        10911 => X"48",  -- 72
        10912 => X"51",  -- 81
        10913 => X"57",  -- 87
        10914 => X"5D",  -- 93
        10915 => X"61",  -- 97
        10916 => X"68",  -- 104
        10917 => X"71",  -- 113
        10918 => X"77",  -- 119
        10919 => X"77",  -- 119
        10920 => X"82",  -- 130
        10921 => X"84",  -- 132
        10922 => X"86",  -- 134
        10923 => X"81",  -- 129
        10924 => X"7B",  -- 123
        10925 => X"78",  -- 120
        10926 => X"7C",  -- 124
        10927 => X"81",  -- 129
        10928 => X"87",  -- 135
        10929 => X"87",  -- 135
        10930 => X"83",  -- 131
        10931 => X"7D",  -- 125
        10932 => X"78",  -- 120
        10933 => X"78",  -- 120
        10934 => X"7D",  -- 125
        10935 => X"81",  -- 129
        10936 => X"8A",  -- 138
        10937 => X"8A",  -- 138
        10938 => X"85",  -- 133
        10939 => X"7D",  -- 125
        10940 => X"79",  -- 121
        10941 => X"7A",  -- 122
        10942 => X"7C",  -- 124
        10943 => X"7E",  -- 126
        10944 => X"7A",  -- 122
        10945 => X"78",  -- 120
        10946 => X"75",  -- 117
        10947 => X"75",  -- 117
        10948 => X"72",  -- 114
        10949 => X"6C",  -- 108
        10950 => X"67",  -- 103
        10951 => X"65",  -- 101
        10952 => X"72",  -- 114
        10953 => X"71",  -- 113
        10954 => X"64",  -- 100
        10955 => X"6D",  -- 109
        10956 => X"58",  -- 88
        10957 => X"65",  -- 101
        10958 => X"4F",  -- 79
        10959 => X"40",  -- 64
        10960 => X"3F",  -- 63
        10961 => X"3C",  -- 60
        10962 => X"3E",  -- 62
        10963 => X"3F",  -- 63
        10964 => X"4A",  -- 74
        10965 => X"4B",  -- 75
        10966 => X"3E",  -- 62
        10967 => X"41",  -- 65
        10968 => X"40",  -- 64
        10969 => X"3F",  -- 63
        10970 => X"27",  -- 39
        10971 => X"2B",  -- 43
        10972 => X"26",  -- 38
        10973 => X"2D",  -- 45
        10974 => X"18",  -- 24
        10975 => X"14",  -- 20
        10976 => X"1D",  -- 29
        10977 => X"22",  -- 34
        10978 => X"1B",  -- 27
        10979 => X"1F",  -- 31
        10980 => X"20",  -- 32
        10981 => X"21",  -- 33
        10982 => X"30",  -- 48
        10983 => X"33",  -- 51
        10984 => X"2E",  -- 46
        10985 => X"29",  -- 41
        10986 => X"23",  -- 35
        10987 => X"23",  -- 35
        10988 => X"26",  -- 38
        10989 => X"29",  -- 41
        10990 => X"29",  -- 41
        10991 => X"25",  -- 37
        10992 => X"27",  -- 39
        10993 => X"24",  -- 36
        10994 => X"26",  -- 38
        10995 => X"2F",  -- 47
        10996 => X"44",  -- 68
        10997 => X"42",  -- 66
        10998 => X"2E",  -- 46
        10999 => X"3A",  -- 58
        11000 => X"4F",  -- 79
        11001 => X"42",  -- 66
        11002 => X"4F",  -- 79
        11003 => X"64",  -- 100
        11004 => X"5A",  -- 90
        11005 => X"58",  -- 88
        11006 => X"4C",  -- 76
        11007 => X"56",  -- 86
        11008 => X"35",  -- 53
        11009 => X"4B",  -- 75
        11010 => X"3F",  -- 63
        11011 => X"2B",  -- 43
        11012 => X"49",  -- 73
        11013 => X"6A",  -- 106
        11014 => X"60",  -- 96
        11015 => X"67",  -- 103
        11016 => X"7D",  -- 125
        11017 => X"75",  -- 117
        11018 => X"7B",  -- 123
        11019 => X"86",  -- 134
        11020 => X"84",  -- 132
        11021 => X"77",  -- 119
        11022 => X"78",  -- 120
        11023 => X"86",  -- 134
        11024 => X"7C",  -- 124
        11025 => X"7D",  -- 125
        11026 => X"7F",  -- 127
        11027 => X"7F",  -- 127
        11028 => X"82",  -- 130
        11029 => X"83",  -- 131
        11030 => X"84",  -- 132
        11031 => X"85",  -- 133
        11032 => X"89",  -- 137
        11033 => X"8D",  -- 141
        11034 => X"8F",  -- 143
        11035 => X"90",  -- 144
        11036 => X"8E",  -- 142
        11037 => X"93",  -- 147
        11038 => X"9E",  -- 158
        11039 => X"A7",  -- 167
        11040 => X"A8",  -- 168
        11041 => X"A5",  -- 165
        11042 => X"A2",  -- 162
        11043 => X"A2",  -- 162
        11044 => X"A4",  -- 164
        11045 => X"AB",  -- 171
        11046 => X"B0",  -- 176
        11047 => X"B3",  -- 179
        11048 => X"A2",  -- 162
        11049 => X"8E",  -- 142
        11050 => X"71",  -- 113
        11051 => X"5D",  -- 93
        11052 => X"58",  -- 88
        11053 => X"5B",  -- 91
        11054 => X"5B",  -- 91
        11055 => X"57",  -- 87
        11056 => X"5C",  -- 92
        11057 => X"5B",  -- 91
        11058 => X"5B",  -- 91
        11059 => X"5E",  -- 94
        11060 => X"66",  -- 102
        11061 => X"6B",  -- 107
        11062 => X"6F",  -- 111
        11063 => X"70",  -- 112
        11064 => X"6A",  -- 106
        11065 => X"69",  -- 105
        11066 => X"69",  -- 105
        11067 => X"69",  -- 105
        11068 => X"6A",  -- 106
        11069 => X"6B",  -- 107
        11070 => X"6B",  -- 107
        11071 => X"6A",  -- 106
        11072 => X"6E",  -- 110
        11073 => X"76",  -- 118
        11074 => X"7A",  -- 122
        11075 => X"74",  -- 116
        11076 => X"6F",  -- 111
        11077 => X"74",  -- 116
        11078 => X"7B",  -- 123
        11079 => X"7E",  -- 126
        11080 => X"77",  -- 119
        11081 => X"78",  -- 120
        11082 => X"7A",  -- 122
        11083 => X"7C",  -- 124
        11084 => X"7C",  -- 124
        11085 => X"7D",  -- 125
        11086 => X"85",  -- 133
        11087 => X"8E",  -- 142
        11088 => X"8A",  -- 138
        11089 => X"8B",  -- 139
        11090 => X"8D",  -- 141
        11091 => X"8B",  -- 139
        11092 => X"89",  -- 137
        11093 => X"8A",  -- 138
        11094 => X"91",  -- 145
        11095 => X"96",  -- 150
        11096 => X"9E",  -- 158
        11097 => X"A4",  -- 164
        11098 => X"A4",  -- 164
        11099 => X"A1",  -- 161
        11100 => X"A4",  -- 164
        11101 => X"AC",  -- 172
        11102 => X"A8",  -- 168
        11103 => X"9D",  -- 157
        11104 => X"A7",  -- 167
        11105 => X"AA",  -- 170
        11106 => X"AC",  -- 172
        11107 => X"A7",  -- 167
        11108 => X"A1",  -- 161
        11109 => X"9F",  -- 159
        11110 => X"9E",  -- 158
        11111 => X"9C",  -- 156
        11112 => X"9E",  -- 158
        11113 => X"A0",  -- 160
        11114 => X"A0",  -- 160
        11115 => X"9F",  -- 159
        11116 => X"9D",  -- 157
        11117 => X"9C",  -- 156
        11118 => X"9E",  -- 158
        11119 => X"A2",  -- 162
        11120 => X"9E",  -- 158
        11121 => X"9F",  -- 159
        11122 => X"9D",  -- 157
        11123 => X"9C",  -- 156
        11124 => X"A0",  -- 160
        11125 => X"A6",  -- 166
        11126 => X"A1",  -- 161
        11127 => X"96",  -- 150
        11128 => X"94",  -- 148
        11129 => X"98",  -- 152
        11130 => X"9D",  -- 157
        11131 => X"A3",  -- 163
        11132 => X"A8",  -- 168
        11133 => X"AB",  -- 171
        11134 => X"AE",  -- 174
        11135 => X"AE",  -- 174
        11136 => X"A8",  -- 168
        11137 => X"AB",  -- 171
        11138 => X"B0",  -- 176
        11139 => X"B1",  -- 177
        11140 => X"AD",  -- 173
        11141 => X"A7",  -- 167
        11142 => X"A2",  -- 162
        11143 => X"9E",  -- 158
        11144 => X"A0",  -- 160
        11145 => X"9C",  -- 156
        11146 => X"99",  -- 153
        11147 => X"9A",  -- 154
        11148 => X"9C",  -- 156
        11149 => X"A0",  -- 160
        11150 => X"A1",  -- 161
        11151 => X"A0",  -- 160
        11152 => X"94",  -- 148
        11153 => X"8A",  -- 138
        11154 => X"7B",  -- 123
        11155 => X"61",  -- 97
        11156 => X"49",  -- 73
        11157 => X"52",  -- 82
        11158 => X"6D",  -- 109
        11159 => X"7C",  -- 124
        11160 => X"95",  -- 149
        11161 => X"9A",  -- 154
        11162 => X"A1",  -- 161
        11163 => X"A0",  -- 160
        11164 => X"9C",  -- 156
        11165 => X"9B",  -- 155
        11166 => X"9E",  -- 158
        11167 => X"A2",  -- 162
        11168 => X"A4",  -- 164
        11169 => X"A4",  -- 164
        11170 => X"9F",  -- 159
        11171 => X"99",  -- 153
        11172 => X"93",  -- 147
        11173 => X"89",  -- 137
        11174 => X"79",  -- 121
        11175 => X"6B",  -- 107
        11176 => X"64",  -- 100
        11177 => X"67",  -- 103
        11178 => X"6D",  -- 109
        11179 => X"78",  -- 120
        11180 => X"89",  -- 137
        11181 => X"9A",  -- 154
        11182 => X"AB",  -- 171
        11183 => X"B4",  -- 180
        11184 => X"AF",  -- 175
        11185 => X"B0",  -- 176
        11186 => X"B0",  -- 176
        11187 => X"B1",  -- 177
        11188 => X"B3",  -- 179
        11189 => X"B3",  -- 179
        11190 => X"B3",  -- 179
        11191 => X"B3",  -- 179
        11192 => X"B3",  -- 179
        11193 => X"BC",  -- 188
        11194 => X"B8",  -- 184
        11195 => X"AE",  -- 174
        11196 => X"B2",  -- 178
        11197 => X"B6",  -- 182
        11198 => X"B4",  -- 180
        11199 => X"B5",  -- 181
        11200 => X"39",  -- 57
        11201 => X"3A",  -- 58
        11202 => X"3B",  -- 59
        11203 => X"3D",  -- 61
        11204 => X"3D",  -- 61
        11205 => X"3F",  -- 63
        11206 => X"40",  -- 64
        11207 => X"40",  -- 64
        11208 => X"3E",  -- 62
        11209 => X"3E",  -- 62
        11210 => X"3F",  -- 63
        11211 => X"40",  -- 64
        11212 => X"40",  -- 64
        11213 => X"40",  -- 64
        11214 => X"40",  -- 64
        11215 => X"40",  -- 64
        11216 => X"41",  -- 65
        11217 => X"41",  -- 65
        11218 => X"41",  -- 65
        11219 => X"40",  -- 64
        11220 => X"3F",  -- 63
        11221 => X"3E",  -- 62
        11222 => X"3C",  -- 60
        11223 => X"3B",  -- 59
        11224 => X"3D",  -- 61
        11225 => X"3F",  -- 63
        11226 => X"44",  -- 68
        11227 => X"47",  -- 71
        11228 => X"4B",  -- 75
        11229 => X"4F",  -- 79
        11230 => X"54",  -- 84
        11231 => X"57",  -- 87
        11232 => X"5C",  -- 92
        11233 => X"64",  -- 100
        11234 => X"6B",  -- 107
        11235 => X"70",  -- 112
        11236 => X"73",  -- 115
        11237 => X"76",  -- 118
        11238 => X"7C",  -- 124
        11239 => X"81",  -- 129
        11240 => X"84",  -- 132
        11241 => X"87",  -- 135
        11242 => X"86",  -- 134
        11243 => X"80",  -- 128
        11244 => X"79",  -- 121
        11245 => X"75",  -- 117
        11246 => X"77",  -- 119
        11247 => X"7B",  -- 123
        11248 => X"7D",  -- 125
        11249 => X"7C",  -- 124
        11250 => X"78",  -- 120
        11251 => X"73",  -- 115
        11252 => X"6F",  -- 111
        11253 => X"72",  -- 114
        11254 => X"76",  -- 118
        11255 => X"7C",  -- 124
        11256 => X"81",  -- 129
        11257 => X"81",  -- 129
        11258 => X"80",  -- 128
        11259 => X"7F",  -- 127
        11260 => X"7F",  -- 127
        11261 => X"7E",  -- 126
        11262 => X"7B",  -- 123
        11263 => X"78",  -- 120
        11264 => X"78",  -- 120
        11265 => X"74",  -- 116
        11266 => X"70",  -- 112
        11267 => X"6F",  -- 111
        11268 => X"6E",  -- 110
        11269 => X"6E",  -- 110
        11270 => X"70",  -- 112
        11271 => X"70",  -- 112
        11272 => X"72",  -- 114
        11273 => X"5F",  -- 95
        11274 => X"48",  -- 72
        11275 => X"48",  -- 72
        11276 => X"32",  -- 50
        11277 => X"38",  -- 56
        11278 => X"2C",  -- 44
        11279 => X"28",  -- 40
        11280 => X"2C",  -- 44
        11281 => X"2F",  -- 47
        11282 => X"31",  -- 49
        11283 => X"39",  -- 57
        11284 => X"49",  -- 73
        11285 => X"4B",  -- 75
        11286 => X"42",  -- 66
        11287 => X"43",  -- 67
        11288 => X"46",  -- 70
        11289 => X"53",  -- 83
        11290 => X"43",  -- 67
        11291 => X"41",  -- 65
        11292 => X"2D",  -- 45
        11293 => X"2B",  -- 43
        11294 => X"13",  -- 19
        11295 => X"10",  -- 16
        11296 => X"22",  -- 34
        11297 => X"1F",  -- 31
        11298 => X"16",  -- 22
        11299 => X"1E",  -- 30
        11300 => X"22",  -- 34
        11301 => X"26",  -- 38
        11302 => X"3D",  -- 61
        11303 => X"48",  -- 72
        11304 => X"43",  -- 67
        11305 => X"48",  -- 72
        11306 => X"46",  -- 70
        11307 => X"3C",  -- 60
        11308 => X"31",  -- 49
        11309 => X"33",  -- 51
        11310 => X"3D",  -- 61
        11311 => X"46",  -- 70
        11312 => X"46",  -- 70
        11313 => X"3D",  -- 61
        11314 => X"35",  -- 53
        11315 => X"38",  -- 56
        11316 => X"41",  -- 65
        11317 => X"35",  -- 53
        11318 => X"25",  -- 37
        11319 => X"2C",  -- 44
        11320 => X"2D",  -- 45
        11321 => X"2A",  -- 42
        11322 => X"38",  -- 56
        11323 => X"42",  -- 66
        11324 => X"4E",  -- 78
        11325 => X"6A",  -- 106
        11326 => X"6D",  -- 109
        11327 => X"6E",  -- 110
        11328 => X"55",  -- 85
        11329 => X"55",  -- 85
        11330 => X"44",  -- 68
        11331 => X"37",  -- 55
        11332 => X"4C",  -- 76
        11333 => X"55",  -- 85
        11334 => X"50",  -- 80
        11335 => X"6D",  -- 109
        11336 => X"7B",  -- 123
        11337 => X"77",  -- 119
        11338 => X"78",  -- 120
        11339 => X"7B",  -- 123
        11340 => X"77",  -- 119
        11341 => X"74",  -- 116
        11342 => X"7B",  -- 123
        11343 => X"89",  -- 137
        11344 => X"77",  -- 119
        11345 => X"7E",  -- 126
        11346 => X"83",  -- 131
        11347 => X"84",  -- 132
        11348 => X"83",  -- 131
        11349 => X"82",  -- 130
        11350 => X"7D",  -- 125
        11351 => X"7A",  -- 122
        11352 => X"87",  -- 135
        11353 => X"90",  -- 144
        11354 => X"9A",  -- 154
        11355 => X"99",  -- 153
        11356 => X"92",  -- 146
        11357 => X"93",  -- 147
        11358 => X"9D",  -- 157
        11359 => X"A9",  -- 169
        11360 => X"AA",  -- 170
        11361 => X"A7",  -- 167
        11362 => X"A4",  -- 164
        11363 => X"A4",  -- 164
        11364 => X"A6",  -- 166
        11365 => X"AA",  -- 170
        11366 => X"B1",  -- 177
        11367 => X"B5",  -- 181
        11368 => X"AB",  -- 171
        11369 => X"A6",  -- 166
        11370 => X"94",  -- 148
        11371 => X"7D",  -- 125
        11372 => X"6F",  -- 111
        11373 => X"66",  -- 102
        11374 => X"59",  -- 89
        11375 => X"4D",  -- 77
        11376 => X"50",  -- 80
        11377 => X"4F",  -- 79
        11378 => X"51",  -- 81
        11379 => X"59",  -- 89
        11380 => X"64",  -- 100
        11381 => X"6E",  -- 110
        11382 => X"72",  -- 114
        11383 => X"73",  -- 115
        11384 => X"6D",  -- 109
        11385 => X"6F",  -- 111
        11386 => X"73",  -- 115
        11387 => X"72",  -- 114
        11388 => X"6F",  -- 111
        11389 => X"6B",  -- 107
        11390 => X"68",  -- 104
        11391 => X"67",  -- 103
        11392 => X"6E",  -- 110
        11393 => X"77",  -- 119
        11394 => X"7B",  -- 123
        11395 => X"76",  -- 118
        11396 => X"75",  -- 117
        11397 => X"7C",  -- 124
        11398 => X"7F",  -- 127
        11399 => X"7C",  -- 124
        11400 => X"76",  -- 118
        11401 => X"76",  -- 118
        11402 => X"79",  -- 121
        11403 => X"7B",  -- 123
        11404 => X"7B",  -- 123
        11405 => X"7C",  -- 124
        11406 => X"83",  -- 131
        11407 => X"8C",  -- 140
        11408 => X"89",  -- 137
        11409 => X"89",  -- 137
        11410 => X"88",  -- 136
        11411 => X"86",  -- 134
        11412 => X"84",  -- 132
        11413 => X"87",  -- 135
        11414 => X"8F",  -- 143
        11415 => X"96",  -- 150
        11416 => X"98",  -- 152
        11417 => X"9A",  -- 154
        11418 => X"98",  -- 152
        11419 => X"98",  -- 152
        11420 => X"9D",  -- 157
        11421 => X"A2",  -- 162
        11422 => X"9F",  -- 159
        11423 => X"96",  -- 150
        11424 => X"9F",  -- 159
        11425 => X"A6",  -- 166
        11426 => X"AB",  -- 171
        11427 => X"A8",  -- 168
        11428 => X"A1",  -- 161
        11429 => X"9F",  -- 159
        11430 => X"9E",  -- 158
        11431 => X"9C",  -- 156
        11432 => X"A0",  -- 160
        11433 => X"A0",  -- 160
        11434 => X"9F",  -- 159
        11435 => X"9D",  -- 157
        11436 => X"9B",  -- 155
        11437 => X"9B",  -- 155
        11438 => X"9D",  -- 157
        11439 => X"A1",  -- 161
        11440 => X"9A",  -- 154
        11441 => X"95",  -- 149
        11442 => X"94",  -- 148
        11443 => X"98",  -- 152
        11444 => X"9E",  -- 158
        11445 => X"9E",  -- 158
        11446 => X"9B",  -- 155
        11447 => X"98",  -- 152
        11448 => X"98",  -- 152
        11449 => X"9B",  -- 155
        11450 => X"9D",  -- 157
        11451 => X"A0",  -- 160
        11452 => X"A3",  -- 163
        11453 => X"A6",  -- 166
        11454 => X"A8",  -- 168
        11455 => X"A9",  -- 169
        11456 => X"A9",  -- 169
        11457 => X"AB",  -- 171
        11458 => X"AF",  -- 175
        11459 => X"AF",  -- 175
        11460 => X"AB",  -- 171
        11461 => X"A4",  -- 164
        11462 => X"9E",  -- 158
        11463 => X"9A",  -- 154
        11464 => X"9F",  -- 159
        11465 => X"9C",  -- 156
        11466 => X"99",  -- 153
        11467 => X"98",  -- 152
        11468 => X"99",  -- 153
        11469 => X"9D",  -- 157
        11470 => X"9E",  -- 158
        11471 => X"9E",  -- 158
        11472 => X"9B",  -- 155
        11473 => X"95",  -- 149
        11474 => X"8A",  -- 138
        11475 => X"6E",  -- 110
        11476 => X"4F",  -- 79
        11477 => X"4D",  -- 77
        11478 => X"65",  -- 101
        11479 => X"75",  -- 117
        11480 => X"8F",  -- 143
        11481 => X"97",  -- 151
        11482 => X"9D",  -- 157
        11483 => X"9D",  -- 157
        11484 => X"99",  -- 153
        11485 => X"9C",  -- 156
        11486 => X"A3",  -- 163
        11487 => X"A7",  -- 167
        11488 => X"A3",  -- 163
        11489 => X"A5",  -- 165
        11490 => X"A4",  -- 164
        11491 => X"A0",  -- 160
        11492 => X"9A",  -- 154
        11493 => X"8D",  -- 141
        11494 => X"79",  -- 121
        11495 => X"69",  -- 105
        11496 => X"63",  -- 99
        11497 => X"61",  -- 97
        11498 => X"63",  -- 99
        11499 => X"70",  -- 112
        11500 => X"86",  -- 134
        11501 => X"9D",  -- 157
        11502 => X"AF",  -- 175
        11503 => X"B7",  -- 183
        11504 => X"B1",  -- 177
        11505 => X"B1",  -- 177
        11506 => X"B0",  -- 176
        11507 => X"B0",  -- 176
        11508 => X"AF",  -- 175
        11509 => X"AE",  -- 174
        11510 => X"AD",  -- 173
        11511 => X"AD",  -- 173
        11512 => X"B0",  -- 176
        11513 => X"BA",  -- 186
        11514 => X"B9",  -- 185
        11515 => X"B4",  -- 180
        11516 => X"B5",  -- 181
        11517 => X"BA",  -- 186
        11518 => X"BB",  -- 187
        11519 => X"BA",  -- 186
        11520 => X"3B",  -- 59
        11521 => X"3B",  -- 59
        11522 => X"3C",  -- 60
        11523 => X"3C",  -- 60
        11524 => X"3E",  -- 62
        11525 => X"3D",  -- 61
        11526 => X"3E",  -- 62
        11527 => X"3F",  -- 63
        11528 => X"40",  -- 64
        11529 => X"40",  -- 64
        11530 => X"40",  -- 64
        11531 => X"41",  -- 65
        11532 => X"40",  -- 64
        11533 => X"41",  -- 65
        11534 => X"41",  -- 65
        11535 => X"41",  -- 65
        11536 => X"41",  -- 65
        11537 => X"3F",  -- 63
        11538 => X"3F",  -- 63
        11539 => X"3E",  -- 62
        11540 => X"3E",  -- 62
        11541 => X"3F",  -- 63
        11542 => X"41",  -- 65
        11543 => X"42",  -- 66
        11544 => X"45",  -- 69
        11545 => X"4B",  -- 75
        11546 => X"51",  -- 81
        11547 => X"58",  -- 88
        11548 => X"5C",  -- 92
        11549 => X"5F",  -- 95
        11550 => X"63",  -- 99
        11551 => X"65",  -- 101
        11552 => X"66",  -- 102
        11553 => X"6B",  -- 107
        11554 => X"72",  -- 114
        11555 => X"76",  -- 118
        11556 => X"76",  -- 118
        11557 => X"77",  -- 119
        11558 => X"7B",  -- 123
        11559 => X"7F",  -- 127
        11560 => X"83",  -- 131
        11561 => X"87",  -- 135
        11562 => X"88",  -- 136
        11563 => X"83",  -- 131
        11564 => X"7B",  -- 123
        11565 => X"74",  -- 116
        11566 => X"74",  -- 116
        11567 => X"77",  -- 119
        11568 => X"73",  -- 115
        11569 => X"73",  -- 115
        11570 => X"72",  -- 114
        11571 => X"70",  -- 112
        11572 => X"6D",  -- 109
        11573 => X"6D",  -- 109
        11574 => X"73",  -- 115
        11575 => X"76",  -- 118
        11576 => X"74",  -- 116
        11577 => X"72",  -- 114
        11578 => X"73",  -- 115
        11579 => X"79",  -- 121
        11580 => X"7D",  -- 125
        11581 => X"7D",  -- 125
        11582 => X"78",  -- 120
        11583 => X"73",  -- 115
        11584 => X"6D",  -- 109
        11585 => X"6E",  -- 110
        11586 => X"72",  -- 114
        11587 => X"73",  -- 115
        11588 => X"74",  -- 116
        11589 => X"70",  -- 112
        11590 => X"6C",  -- 108
        11591 => X"67",  -- 103
        11592 => X"51",  -- 81
        11593 => X"3C",  -- 60
        11594 => X"2B",  -- 43
        11595 => X"2F",  -- 47
        11596 => X"23",  -- 35
        11597 => X"26",  -- 38
        11598 => X"2C",  -- 44
        11599 => X"39",  -- 57
        11600 => X"2D",  -- 45
        11601 => X"34",  -- 52
        11602 => X"33",  -- 51
        11603 => X"3D",  -- 61
        11604 => X"4E",  -- 78
        11605 => X"51",  -- 81
        11606 => X"4F",  -- 79
        11607 => X"4E",  -- 78
        11608 => X"45",  -- 69
        11609 => X"65",  -- 101
        11610 => X"6C",  -- 108
        11611 => X"60",  -- 96
        11612 => X"41",  -- 65
        11613 => X"32",  -- 50
        11614 => X"22",  -- 34
        11615 => X"25",  -- 37
        11616 => X"1C",  -- 28
        11617 => X"20",  -- 32
        11618 => X"1F",  -- 31
        11619 => X"2F",  -- 47
        11620 => X"37",  -- 55
        11621 => X"39",  -- 57
        11622 => X"52",  -- 82
        11623 => X"61",  -- 97
        11624 => X"55",  -- 85
        11625 => X"60",  -- 96
        11626 => X"66",  -- 102
        11627 => X"5E",  -- 94
        11628 => X"56",  -- 86
        11629 => X"5B",  -- 91
        11630 => X"69",  -- 105
        11631 => X"76",  -- 118
        11632 => X"7C",  -- 124
        11633 => X"71",  -- 113
        11634 => X"5D",  -- 93
        11635 => X"56",  -- 86
        11636 => X"51",  -- 81
        11637 => X"43",  -- 67
        11638 => X"42",  -- 66
        11639 => X"49",  -- 73
        11640 => X"30",  -- 48
        11641 => X"25",  -- 37
        11642 => X"2A",  -- 42
        11643 => X"28",  -- 40
        11644 => X"39",  -- 57
        11645 => X"5B",  -- 91
        11646 => X"6E",  -- 110
        11647 => X"74",  -- 116
        11648 => X"76",  -- 118
        11649 => X"5E",  -- 94
        11650 => X"55",  -- 85
        11651 => X"4A",  -- 74
        11652 => X"41",  -- 65
        11653 => X"41",  -- 65
        11654 => X"4F",  -- 79
        11655 => X"71",  -- 113
        11656 => X"66",  -- 102
        11657 => X"6F",  -- 111
        11658 => X"77",  -- 119
        11659 => X"77",  -- 119
        11660 => X"76",  -- 118
        11661 => X"79",  -- 121
        11662 => X"7C",  -- 124
        11663 => X"80",  -- 128
        11664 => X"7C",  -- 124
        11665 => X"82",  -- 130
        11666 => X"85",  -- 133
        11667 => X"83",  -- 131
        11668 => X"83",  -- 131
        11669 => X"84",  -- 132
        11670 => X"82",  -- 130
        11671 => X"7F",  -- 127
        11672 => X"85",  -- 133
        11673 => X"86",  -- 134
        11674 => X"8B",  -- 139
        11675 => X"92",  -- 146
        11676 => X"9A",  -- 154
        11677 => X"9F",  -- 159
        11678 => X"9E",  -- 158
        11679 => X"9D",  -- 157
        11680 => X"AC",  -- 172
        11681 => X"AD",  -- 173
        11682 => X"AD",  -- 173
        11683 => X"AB",  -- 171
        11684 => X"A9",  -- 169
        11685 => X"AA",  -- 170
        11686 => X"AE",  -- 174
        11687 => X"B2",  -- 178
        11688 => X"AF",  -- 175
        11689 => X"AD",  -- 173
        11690 => X"9B",  -- 155
        11691 => X"7C",  -- 124
        11692 => X"64",  -- 100
        11693 => X"5C",  -- 92
        11694 => X"59",  -- 89
        11695 => X"57",  -- 87
        11696 => X"56",  -- 86
        11697 => X"54",  -- 84
        11698 => X"55",  -- 85
        11699 => X"5B",  -- 91
        11700 => X"64",  -- 100
        11701 => X"6A",  -- 106
        11702 => X"6A",  -- 106
        11703 => X"6A",  -- 106
        11704 => X"79",  -- 121
        11705 => X"7B",  -- 123
        11706 => X"78",  -- 120
        11707 => X"71",  -- 113
        11708 => X"68",  -- 104
        11709 => X"66",  -- 102
        11710 => X"6B",  -- 107
        11711 => X"72",  -- 114
        11712 => X"75",  -- 117
        11713 => X"79",  -- 121
        11714 => X"7D",  -- 125
        11715 => X"7C",  -- 124
        11716 => X"80",  -- 128
        11717 => X"84",  -- 132
        11718 => X"80",  -- 128
        11719 => X"77",  -- 119
        11720 => X"75",  -- 117
        11721 => X"71",  -- 113
        11722 => X"71",  -- 113
        11723 => X"75",  -- 117
        11724 => X"7B",  -- 123
        11725 => X"7D",  -- 125
        11726 => X"80",  -- 128
        11727 => X"85",  -- 133
        11728 => X"88",  -- 136
        11729 => X"86",  -- 134
        11730 => X"83",  -- 131
        11731 => X"7E",  -- 126
        11732 => X"7D",  -- 125
        11733 => X"82",  -- 130
        11734 => X"8D",  -- 141
        11735 => X"96",  -- 150
        11736 => X"96",  -- 150
        11737 => X"92",  -- 146
        11738 => X"91",  -- 145
        11739 => X"97",  -- 151
        11740 => X"9A",  -- 154
        11741 => X"97",  -- 151
        11742 => X"96",  -- 150
        11743 => X"99",  -- 153
        11744 => X"97",  -- 151
        11745 => X"A1",  -- 161
        11746 => X"A8",  -- 168
        11747 => X"A7",  -- 167
        11748 => X"A4",  -- 164
        11749 => X"A1",  -- 161
        11750 => X"9D",  -- 157
        11751 => X"9A",  -- 154
        11752 => X"A1",  -- 161
        11753 => X"A0",  -- 160
        11754 => X"9E",  -- 158
        11755 => X"9C",  -- 156
        11756 => X"9B",  -- 155
        11757 => X"9D",  -- 157
        11758 => X"9F",  -- 159
        11759 => X"A2",  -- 162
        11760 => X"9E",  -- 158
        11761 => X"92",  -- 146
        11762 => X"8F",  -- 143
        11763 => X"96",  -- 150
        11764 => X"96",  -- 150
        11765 => X"8E",  -- 142
        11766 => X"90",  -- 144
        11767 => X"9B",  -- 155
        11768 => X"A0",  -- 160
        11769 => X"9F",  -- 159
        11770 => X"9F",  -- 159
        11771 => X"9F",  -- 159
        11772 => X"A1",  -- 161
        11773 => X"A4",  -- 164
        11774 => X"A6",  -- 166
        11775 => X"A8",  -- 168
        11776 => X"AA",  -- 170
        11777 => X"AB",  -- 171
        11778 => X"AD",  -- 173
        11779 => X"AD",  -- 173
        11780 => X"AA",  -- 170
        11781 => X"A6",  -- 166
        11782 => X"A1",  -- 161
        11783 => X"9D",  -- 157
        11784 => X"A3",  -- 163
        11785 => X"A0",  -- 160
        11786 => X"9C",  -- 156
        11787 => X"9A",  -- 154
        11788 => X"99",  -- 153
        11789 => X"9B",  -- 155
        11790 => X"9C",  -- 156
        11791 => X"9D",  -- 157
        11792 => X"A5",  -- 165
        11793 => X"9A",  -- 154
        11794 => X"90",  -- 144
        11795 => X"7A",  -- 122
        11796 => X"59",  -- 89
        11797 => X"49",  -- 73
        11798 => X"59",  -- 89
        11799 => X"6A",  -- 106
        11800 => X"7B",  -- 123
        11801 => X"8A",  -- 138
        11802 => X"9A",  -- 154
        11803 => X"9F",  -- 159
        11804 => X"9F",  -- 159
        11805 => X"A2",  -- 162
        11806 => X"A6",  -- 166
        11807 => X"A8",  -- 168
        11808 => X"A2",  -- 162
        11809 => X"A5",  -- 165
        11810 => X"A7",  -- 167
        11811 => X"A5",  -- 165
        11812 => X"A2",  -- 162
        11813 => X"98",  -- 152
        11814 => X"86",  -- 134
        11815 => X"77",  -- 119
        11816 => X"6B",  -- 107
        11817 => X"62",  -- 98
        11818 => X"5D",  -- 93
        11819 => X"6B",  -- 107
        11820 => X"88",  -- 136
        11821 => X"A3",  -- 163
        11822 => X"B2",  -- 178
        11823 => X"B6",  -- 182
        11824 => X"B3",  -- 179
        11825 => X"B1",  -- 177
        11826 => X"B0",  -- 176
        11827 => X"AF",  -- 175
        11828 => X"AF",  -- 175
        11829 => X"AF",  -- 175
        11830 => X"AF",  -- 175
        11831 => X"AE",  -- 174
        11832 => X"B5",  -- 181
        11833 => X"B9",  -- 185
        11834 => X"BC",  -- 188
        11835 => X"BA",  -- 186
        11836 => X"B6",  -- 182
        11837 => X"BA",  -- 186
        11838 => X"BA",  -- 186
        11839 => X"B4",  -- 180
        11840 => X"3A",  -- 58
        11841 => X"3A",  -- 58
        11842 => X"3C",  -- 60
        11843 => X"3C",  -- 60
        11844 => X"3D",  -- 61
        11845 => X"3D",  -- 61
        11846 => X"3E",  -- 62
        11847 => X"3E",  -- 62
        11848 => X"3F",  -- 63
        11849 => X"3F",  -- 63
        11850 => X"3E",  -- 62
        11851 => X"3D",  -- 61
        11852 => X"3C",  -- 60
        11853 => X"3D",  -- 61
        11854 => X"3E",  -- 62
        11855 => X"3E",  -- 62
        11856 => X"3F",  -- 63
        11857 => X"3F",  -- 63
        11858 => X"3F",  -- 63
        11859 => X"42",  -- 66
        11860 => X"45",  -- 69
        11861 => X"49",  -- 73
        11862 => X"4F",  -- 79
        11863 => X"51",  -- 81
        11864 => X"55",  -- 85
        11865 => X"5B",  -- 91
        11866 => X"63",  -- 99
        11867 => X"68",  -- 104
        11868 => X"6B",  -- 107
        11869 => X"6B",  -- 107
        11870 => X"6D",  -- 109
        11871 => X"6E",  -- 110
        11872 => X"6D",  -- 109
        11873 => X"6F",  -- 111
        11874 => X"72",  -- 114
        11875 => X"74",  -- 116
        11876 => X"73",  -- 115
        11877 => X"70",  -- 112
        11878 => X"73",  -- 115
        11879 => X"79",  -- 121
        11880 => X"7F",  -- 127
        11881 => X"83",  -- 131
        11882 => X"85",  -- 133
        11883 => X"82",  -- 130
        11884 => X"79",  -- 121
        11885 => X"74",  -- 116
        11886 => X"74",  -- 116
        11887 => X"76",  -- 118
        11888 => X"75",  -- 117
        11889 => X"76",  -- 118
        11890 => X"77",  -- 119
        11891 => X"76",  -- 118
        11892 => X"73",  -- 115
        11893 => X"72",  -- 114
        11894 => X"74",  -- 116
        11895 => X"77",  -- 119
        11896 => X"71",  -- 113
        11897 => X"6E",  -- 110
        11898 => X"6C",  -- 108
        11899 => X"71",  -- 113
        11900 => X"77",  -- 119
        11901 => X"76",  -- 118
        11902 => X"73",  -- 115
        11903 => X"70",  -- 112
        11904 => X"63",  -- 99
        11905 => X"6D",  -- 109
        11906 => X"75",  -- 117
        11907 => X"78",  -- 120
        11908 => X"72",  -- 114
        11909 => X"64",  -- 100
        11910 => X"52",  -- 82
        11911 => X"43",  -- 67
        11912 => X"38",  -- 56
        11913 => X"25",  -- 37
        11914 => X"1F",  -- 31
        11915 => X"25",  -- 37
        11916 => X"21",  -- 33
        11917 => X"30",  -- 48
        11918 => X"4F",  -- 79
        11919 => X"6A",  -- 106
        11920 => X"52",  -- 82
        11921 => X"5E",  -- 94
        11922 => X"58",  -- 88
        11923 => X"61",  -- 97
        11924 => X"6C",  -- 108
        11925 => X"6E",  -- 110
        11926 => X"71",  -- 113
        11927 => X"6C",  -- 108
        11928 => X"66",  -- 102
        11929 => X"77",  -- 119
        11930 => X"78",  -- 120
        11931 => X"69",  -- 105
        11932 => X"64",  -- 100
        11933 => X"55",  -- 85
        11934 => X"3F",  -- 63
        11935 => X"2D",  -- 45
        11936 => X"1C",  -- 28
        11937 => X"2A",  -- 42
        11938 => X"37",  -- 55
        11939 => X"4D",  -- 77
        11940 => X"57",  -- 87
        11941 => X"58",  -- 88
        11942 => X"6E",  -- 110
        11943 => X"78",  -- 120
        11944 => X"6E",  -- 110
        11945 => X"76",  -- 118
        11946 => X"78",  -- 120
        11947 => X"7A",  -- 122
        11948 => X"7E",  -- 126
        11949 => X"89",  -- 137
        11950 => X"8C",  -- 140
        11951 => X"89",  -- 137
        11952 => X"8D",  -- 141
        11953 => X"8E",  -- 142
        11954 => X"85",  -- 133
        11955 => X"85",  -- 133
        11956 => X"7B",  -- 123
        11957 => X"69",  -- 105
        11958 => X"6B",  -- 107
        11959 => X"66",  -- 102
        11960 => X"4D",  -- 77
        11961 => X"2E",  -- 46
        11962 => X"2D",  -- 45
        11963 => X"22",  -- 34
        11964 => X"28",  -- 40
        11965 => X"33",  -- 51
        11966 => X"4C",  -- 76
        11967 => X"61",  -- 97
        11968 => X"6E",  -- 110
        11969 => X"66",  -- 102
        11970 => X"74",  -- 116
        11971 => X"64",  -- 100
        11972 => X"48",  -- 72
        11973 => X"4A",  -- 74
        11974 => X"51",  -- 81
        11975 => X"57",  -- 87
        11976 => X"5E",  -- 94
        11977 => X"69",  -- 105
        11978 => X"70",  -- 112
        11979 => X"6F",  -- 111
        11980 => X"71",  -- 113
        11981 => X"7C",  -- 124
        11982 => X"81",  -- 129
        11983 => X"80",  -- 128
        11984 => X"7C",  -- 124
        11985 => X"80",  -- 128
        11986 => X"7F",  -- 127
        11987 => X"78",  -- 120
        11988 => X"78",  -- 120
        11989 => X"82",  -- 130
        11990 => X"88",  -- 136
        11991 => X"8A",  -- 138
        11992 => X"84",  -- 132
        11993 => X"89",  -- 137
        11994 => X"90",  -- 144
        11995 => X"97",  -- 151
        11996 => X"9D",  -- 157
        11997 => X"9D",  -- 157
        11998 => X"9C",  -- 156
        11999 => X"9A",  -- 154
        12000 => X"A9",  -- 169
        12001 => X"AD",  -- 173
        12002 => X"B2",  -- 178
        12003 => X"B0",  -- 176
        12004 => X"AC",  -- 172
        12005 => X"AA",  -- 170
        12006 => X"A9",  -- 169
        12007 => X"AC",  -- 172
        12008 => X"AD",  -- 173
        12009 => X"A9",  -- 169
        12010 => X"97",  -- 151
        12011 => X"7A",  -- 122
        12012 => X"5E",  -- 94
        12013 => X"50",  -- 80
        12014 => X"51",  -- 81
        12015 => X"53",  -- 83
        12016 => X"61",  -- 97
        12017 => X"5E",  -- 94
        12018 => X"5E",  -- 94
        12019 => X"61",  -- 97
        12020 => X"65",  -- 101
        12021 => X"6A",  -- 106
        12022 => X"6B",  -- 107
        12023 => X"69",  -- 105
        12024 => X"76",  -- 118
        12025 => X"7A",  -- 122
        12026 => X"7B",  -- 123
        12027 => X"76",  -- 118
        12028 => X"6E",  -- 110
        12029 => X"6A",  -- 106
        12030 => X"6D",  -- 109
        12031 => X"71",  -- 113
        12032 => X"79",  -- 121
        12033 => X"77",  -- 119
        12034 => X"78",  -- 120
        12035 => X"7D",  -- 125
        12036 => X"82",  -- 130
        12037 => X"80",  -- 128
        12038 => X"76",  -- 118
        12039 => X"6D",  -- 109
        12040 => X"72",  -- 114
        12041 => X"6C",  -- 108
        12042 => X"69",  -- 105
        12043 => X"70",  -- 112
        12044 => X"79",  -- 121
        12045 => X"7D",  -- 125
        12046 => X"7E",  -- 126
        12047 => X"7F",  -- 127
        12048 => X"85",  -- 133
        12049 => X"82",  -- 130
        12050 => X"7E",  -- 126
        12051 => X"79",  -- 121
        12052 => X"78",  -- 120
        12053 => X"7D",  -- 125
        12054 => X"8A",  -- 138
        12055 => X"94",  -- 148
        12056 => X"96",  -- 150
        12057 => X"90",  -- 144
        12058 => X"91",  -- 145
        12059 => X"98",  -- 152
        12060 => X"99",  -- 153
        12061 => X"93",  -- 147
        12062 => X"95",  -- 149
        12063 => X"9D",  -- 157
        12064 => X"95",  -- 149
        12065 => X"9D",  -- 157
        12066 => X"A5",  -- 165
        12067 => X"A5",  -- 165
        12068 => X"A4",  -- 164
        12069 => X"A1",  -- 161
        12070 => X"9D",  -- 157
        12071 => X"98",  -- 152
        12072 => X"A1",  -- 161
        12073 => X"A0",  -- 160
        12074 => X"9E",  -- 158
        12075 => X"9C",  -- 156
        12076 => X"9C",  -- 156
        12077 => X"9E",  -- 158
        12078 => X"A0",  -- 160
        12079 => X"A2",  -- 162
        12080 => X"A1",  -- 161
        12081 => X"95",  -- 149
        12082 => X"90",  -- 144
        12083 => X"91",  -- 145
        12084 => X"8B",  -- 139
        12085 => X"84",  -- 132
        12086 => X"8C",  -- 140
        12087 => X"9C",  -- 156
        12088 => X"A0",  -- 160
        12089 => X"9F",  -- 159
        12090 => X"9F",  -- 159
        12091 => X"A0",  -- 160
        12092 => X"A3",  -- 163
        12093 => X"A6",  -- 166
        12094 => X"A9",  -- 169
        12095 => X"AC",  -- 172
        12096 => X"A9",  -- 169
        12097 => X"AB",  -- 171
        12098 => X"AC",  -- 172
        12099 => X"AE",  -- 174
        12100 => X"AE",  -- 174
        12101 => X"AC",  -- 172
        12102 => X"A8",  -- 168
        12103 => X"A5",  -- 165
        12104 => X"A1",  -- 161
        12105 => X"9F",  -- 159
        12106 => X"9B",  -- 155
        12107 => X"98",  -- 152
        12108 => X"96",  -- 150
        12109 => X"96",  -- 150
        12110 => X"98",  -- 152
        12111 => X"99",  -- 153
        12112 => X"A8",  -- 168
        12113 => X"9B",  -- 155
        12114 => X"92",  -- 146
        12115 => X"80",  -- 128
        12116 => X"5D",  -- 93
        12117 => X"45",  -- 69
        12118 => X"4B",  -- 75
        12119 => X"56",  -- 86
        12120 => X"5F",  -- 95
        12121 => X"79",  -- 121
        12122 => X"95",  -- 149
        12123 => X"A1",  -- 161
        12124 => X"A5",  -- 165
        12125 => X"A7",  -- 167
        12126 => X"A5",  -- 165
        12127 => X"A2",  -- 162
        12128 => X"A1",  -- 161
        12129 => X"A3",  -- 163
        12130 => X"A4",  -- 164
        12131 => X"A3",  -- 163
        12132 => X"A5",  -- 165
        12133 => X"A2",  -- 162
        12134 => X"96",  -- 150
        12135 => X"8B",  -- 139
        12136 => X"76",  -- 118
        12137 => X"68",  -- 104
        12138 => X"60",  -- 96
        12139 => X"6D",  -- 109
        12140 => X"8D",  -- 141
        12141 => X"A7",  -- 167
        12142 => X"B4",  -- 180
        12143 => X"B3",  -- 179
        12144 => X"B3",  -- 179
        12145 => X"B2",  -- 178
        12146 => X"B0",  -- 176
        12147 => X"B0",  -- 176
        12148 => X"B2",  -- 178
        12149 => X"B4",  -- 180
        12150 => X"B7",  -- 183
        12151 => X"BA",  -- 186
        12152 => X"BA",  -- 186
        12153 => X"BC",  -- 188
        12154 => X"BF",  -- 191
        12155 => X"BE",  -- 190
        12156 => X"B7",  -- 183
        12157 => X"B9",  -- 185
        12158 => X"B6",  -- 182
        12159 => X"A6",  -- 166
        12160 => X"3A",  -- 58
        12161 => X"3A",  -- 58
        12162 => X"3C",  -- 60
        12163 => X"3C",  -- 60
        12164 => X"3C",  -- 60
        12165 => X"3C",  -- 60
        12166 => X"3D",  -- 61
        12167 => X"3E",  -- 62
        12168 => X"3C",  -- 60
        12169 => X"3C",  -- 60
        12170 => X"3D",  -- 61
        12171 => X"3E",  -- 62
        12172 => X"3E",  -- 62
        12173 => X"40",  -- 64
        12174 => X"42",  -- 66
        12175 => X"44",  -- 68
        12176 => X"4B",  -- 75
        12177 => X"4C",  -- 76
        12178 => X"50",  -- 80
        12179 => X"54",  -- 84
        12180 => X"59",  -- 89
        12181 => X"5F",  -- 95
        12182 => X"64",  -- 100
        12183 => X"66",  -- 102
        12184 => X"67",  -- 103
        12185 => X"6C",  -- 108
        12186 => X"6F",  -- 111
        12187 => X"70",  -- 112
        12188 => X"6E",  -- 110
        12189 => X"6B",  -- 107
        12190 => X"6B",  -- 107
        12191 => X"6D",  -- 109
        12192 => X"6B",  -- 107
        12193 => X"6A",  -- 106
        12194 => X"6B",  -- 107
        12195 => X"6D",  -- 109
        12196 => X"6B",  -- 107
        12197 => X"67",  -- 103
        12198 => X"69",  -- 105
        12199 => X"6E",  -- 110
        12200 => X"77",  -- 119
        12201 => X"7C",  -- 124
        12202 => X"81",  -- 129
        12203 => X"80",  -- 128
        12204 => X"7C",  -- 124
        12205 => X"7B",  -- 123
        12206 => X"7F",  -- 127
        12207 => X"82",  -- 130
        12208 => X"87",  -- 135
        12209 => X"89",  -- 137
        12210 => X"88",  -- 136
        12211 => X"83",  -- 131
        12212 => X"7D",  -- 125
        12213 => X"7A",  -- 122
        12214 => X"7A",  -- 122
        12215 => X"7B",  -- 123
        12216 => X"79",  -- 121
        12217 => X"72",  -- 114
        12218 => X"6E",  -- 110
        12219 => X"6F",  -- 111
        12220 => X"70",  -- 112
        12221 => X"6D",  -- 109
        12222 => X"6B",  -- 107
        12223 => X"6C",  -- 108
        12224 => X"70",  -- 112
        12225 => X"73",  -- 115
        12226 => X"72",  -- 114
        12227 => X"68",  -- 104
        12228 => X"5A",  -- 90
        12229 => X"4A",  -- 74
        12230 => X"37",  -- 55
        12231 => X"27",  -- 39
        12232 => X"21",  -- 33
        12233 => X"1F",  -- 31
        12234 => X"23",  -- 35
        12235 => X"25",  -- 37
        12236 => X"2A",  -- 42
        12237 => X"43",  -- 67
        12238 => X"68",  -- 104
        12239 => X"7C",  -- 124
        12240 => X"7C",  -- 124
        12241 => X"8C",  -- 140
        12242 => X"82",  -- 130
        12243 => X"86",  -- 134
        12244 => X"8C",  -- 140
        12245 => X"84",  -- 132
        12246 => X"89",  -- 137
        12247 => X"83",  -- 131
        12248 => X"7E",  -- 126
        12249 => X"74",  -- 116
        12250 => X"66",  -- 102
        12251 => X"51",  -- 81
        12252 => X"6F",  -- 111
        12253 => X"6A",  -- 106
        12254 => X"55",  -- 85
        12255 => X"2E",  -- 46
        12256 => X"20",  -- 32
        12257 => X"37",  -- 55
        12258 => X"47",  -- 71
        12259 => X"5A",  -- 90
        12260 => X"5C",  -- 92
        12261 => X"5C",  -- 92
        12262 => X"6E",  -- 110
        12263 => X"76",  -- 118
        12264 => X"77",  -- 119
        12265 => X"76",  -- 118
        12266 => X"72",  -- 114
        12267 => X"73",  -- 115
        12268 => X"7E",  -- 126
        12269 => X"8C",  -- 140
        12270 => X"8C",  -- 140
        12271 => X"81",  -- 129
        12272 => X"82",  -- 130
        12273 => X"90",  -- 144
        12274 => X"94",  -- 148
        12275 => X"9C",  -- 156
        12276 => X"94",  -- 148
        12277 => X"85",  -- 133
        12278 => X"86",  -- 134
        12279 => X"73",  -- 115
        12280 => X"6A",  -- 106
        12281 => X"4F",  -- 79
        12282 => X"4A",  -- 74
        12283 => X"2F",  -- 47
        12284 => X"22",  -- 34
        12285 => X"1C",  -- 28
        12286 => X"2F",  -- 47
        12287 => X"43",  -- 67
        12288 => X"4F",  -- 79
        12289 => X"5C",  -- 92
        12290 => X"78",  -- 120
        12291 => X"71",  -- 113
        12292 => X"63",  -- 99
        12293 => X"69",  -- 105
        12294 => X"5F",  -- 95
        12295 => X"54",  -- 84
        12296 => X"5E",  -- 94
        12297 => X"64",  -- 100
        12298 => X"69",  -- 105
        12299 => X"6D",  -- 109
        12300 => X"73",  -- 115
        12301 => X"7B",  -- 123
        12302 => X"82",  -- 130
        12303 => X"85",  -- 133
        12304 => X"7B",  -- 123
        12305 => X"80",  -- 128
        12306 => X"7D",  -- 125
        12307 => X"75",  -- 117
        12308 => X"74",  -- 116
        12309 => X"80",  -- 128
        12310 => X"8A",  -- 138
        12311 => X"8D",  -- 141
        12312 => X"85",  -- 133
        12313 => X"90",  -- 144
        12314 => X"9A",  -- 154
        12315 => X"9F",  -- 159
        12316 => X"9E",  -- 158
        12317 => X"9C",  -- 156
        12318 => X"9F",  -- 159
        12319 => X"A1",  -- 161
        12320 => X"A6",  -- 166
        12321 => X"AC",  -- 172
        12322 => X"B3",  -- 179
        12323 => X"B5",  -- 181
        12324 => X"B0",  -- 176
        12325 => X"AB",  -- 171
        12326 => X"AB",  -- 171
        12327 => X"AC",  -- 172
        12328 => X"B6",  -- 182
        12329 => X"B0",  -- 176
        12330 => X"A6",  -- 166
        12331 => X"97",  -- 151
        12332 => X"83",  -- 131
        12333 => X"6E",  -- 110
        12334 => X"5E",  -- 94
        12335 => X"58",  -- 88
        12336 => X"60",  -- 96
        12337 => X"5F",  -- 95
        12338 => X"5E",  -- 94
        12339 => X"60",  -- 96
        12340 => X"63",  -- 99
        12341 => X"6A",  -- 106
        12342 => X"70",  -- 112
        12343 => X"74",  -- 116
        12344 => X"70",  -- 112
        12345 => X"73",  -- 115
        12346 => X"79",  -- 121
        12347 => X"7B",  -- 123
        12348 => X"7B",  -- 123
        12349 => X"77",  -- 119
        12350 => X"73",  -- 115
        12351 => X"70",  -- 112
        12352 => X"79",  -- 121
        12353 => X"73",  -- 115
        12354 => X"75",  -- 117
        12355 => X"7D",  -- 125
        12356 => X"80",  -- 128
        12357 => X"78",  -- 120
        12358 => X"6F",  -- 111
        12359 => X"6C",  -- 108
        12360 => X"70",  -- 112
        12361 => X"6A",  -- 106
        12362 => X"69",  -- 105
        12363 => X"70",  -- 112
        12364 => X"7A",  -- 122
        12365 => X"7E",  -- 126
        12366 => X"7F",  -- 127
        12367 => X"7F",  -- 127
        12368 => X"81",  -- 129
        12369 => X"80",  -- 128
        12370 => X"7E",  -- 126
        12371 => X"7A",  -- 122
        12372 => X"78",  -- 120
        12373 => X"7D",  -- 125
        12374 => X"88",  -- 136
        12375 => X"91",  -- 145
        12376 => X"94",  -- 148
        12377 => X"93",  -- 147
        12378 => X"92",  -- 146
        12379 => X"94",  -- 148
        12380 => X"96",  -- 150
        12381 => X"96",  -- 150
        12382 => X"98",  -- 152
        12383 => X"9B",  -- 155
        12384 => X"97",  -- 151
        12385 => X"9C",  -- 156
        12386 => X"A1",  -- 161
        12387 => X"A2",  -- 162
        12388 => X"A2",  -- 162
        12389 => X"A2",  -- 162
        12390 => X"9E",  -- 158
        12391 => X"98",  -- 152
        12392 => X"9D",  -- 157
        12393 => X"9C",  -- 156
        12394 => X"99",  -- 153
        12395 => X"99",  -- 153
        12396 => X"9A",  -- 154
        12397 => X"9C",  -- 156
        12398 => X"9D",  -- 157
        12399 => X"9E",  -- 158
        12400 => X"97",  -- 151
        12401 => X"95",  -- 149
        12402 => X"8E",  -- 142
        12403 => X"85",  -- 133
        12404 => X"80",  -- 128
        12405 => X"85",  -- 133
        12406 => X"90",  -- 144
        12407 => X"98",  -- 152
        12408 => X"99",  -- 153
        12409 => X"9B",  -- 155
        12410 => X"9D",  -- 157
        12411 => X"A1",  -- 161
        12412 => X"A4",  -- 164
        12413 => X"A7",  -- 167
        12414 => X"A9",  -- 169
        12415 => X"AA",  -- 170
        12416 => X"A7",  -- 167
        12417 => X"A8",  -- 168
        12418 => X"AD",  -- 173
        12419 => X"B1",  -- 177
        12420 => X"B2",  -- 178
        12421 => X"B0",  -- 176
        12422 => X"AB",  -- 171
        12423 => X"A6",  -- 166
        12424 => X"9D",  -- 157
        12425 => X"9C",  -- 156
        12426 => X"99",  -- 153
        12427 => X"95",  -- 149
        12428 => X"93",  -- 147
        12429 => X"93",  -- 147
        12430 => X"96",  -- 150
        12431 => X"97",  -- 151
        12432 => X"9F",  -- 159
        12433 => X"9A",  -- 154
        12434 => X"95",  -- 149
        12435 => X"7E",  -- 126
        12436 => X"57",  -- 87
        12437 => X"43",  -- 67
        12438 => X"42",  -- 66
        12439 => X"44",  -- 68
        12440 => X"4A",  -- 74
        12441 => X"68",  -- 104
        12442 => X"8A",  -- 138
        12443 => X"9B",  -- 155
        12444 => X"A2",  -- 162
        12445 => X"A5",  -- 165
        12446 => X"A2",  -- 162
        12447 => X"9E",  -- 158
        12448 => X"9C",  -- 156
        12449 => X"9F",  -- 159
        12450 => X"A2",  -- 162
        12451 => X"A4",  -- 164
        12452 => X"A6",  -- 166
        12453 => X"A4",  -- 164
        12454 => X"99",  -- 153
        12455 => X"8E",  -- 142
        12456 => X"76",  -- 118
        12457 => X"6A",  -- 106
        12458 => X"62",  -- 98
        12459 => X"6F",  -- 111
        12460 => X"8D",  -- 141
        12461 => X"A6",  -- 166
        12462 => X"B2",  -- 178
        12463 => X"B1",  -- 177
        12464 => X"B3",  -- 179
        12465 => X"B2",  -- 178
        12466 => X"B0",  -- 176
        12467 => X"B0",  -- 176
        12468 => X"B2",  -- 178
        12469 => X"B8",  -- 184
        12470 => X"BE",  -- 190
        12471 => X"C0",  -- 192
        12472 => X"C0",  -- 192
        12473 => X"BC",  -- 188
        12474 => X"C2",  -- 194
        12475 => X"C0",  -- 192
        12476 => X"B8",  -- 184
        12477 => X"BA",  -- 186
        12478 => X"B4",  -- 180
        12479 => X"9F",  -- 159
        12480 => X"3A",  -- 58
        12481 => X"3B",  -- 59
        12482 => X"3A",  -- 58
        12483 => X"3B",  -- 59
        12484 => X"3C",  -- 60
        12485 => X"3D",  -- 61
        12486 => X"3D",  -- 61
        12487 => X"3E",  -- 62
        12488 => X"3E",  -- 62
        12489 => X"3E",  -- 62
        12490 => X"40",  -- 64
        12491 => X"44",  -- 68
        12492 => X"47",  -- 71
        12493 => X"4C",  -- 76
        12494 => X"50",  -- 80
        12495 => X"52",  -- 82
        12496 => X"59",  -- 89
        12497 => X"5C",  -- 92
        12498 => X"61",  -- 97
        12499 => X"67",  -- 103
        12500 => X"6E",  -- 110
        12501 => X"73",  -- 115
        12502 => X"75",  -- 117
        12503 => X"77",  -- 119
        12504 => X"72",  -- 114
        12505 => X"75",  -- 117
        12506 => X"75",  -- 117
        12507 => X"71",  -- 113
        12508 => X"6A",  -- 106
        12509 => X"64",  -- 100
        12510 => X"64",  -- 100
        12511 => X"65",  -- 101
        12512 => X"69",  -- 105
        12513 => X"65",  -- 101
        12514 => X"63",  -- 99
        12515 => X"65",  -- 101
        12516 => X"64",  -- 100
        12517 => X"60",  -- 96
        12518 => X"62",  -- 98
        12519 => X"66",  -- 102
        12520 => X"75",  -- 117
        12521 => X"7B",  -- 123
        12522 => X"81",  -- 129
        12523 => X"82",  -- 130
        12524 => X"83",  -- 131
        12525 => X"87",  -- 135
        12526 => X"8F",  -- 143
        12527 => X"97",  -- 151
        12528 => X"99",  -- 153
        12529 => X"98",  -- 152
        12530 => X"96",  -- 150
        12531 => X"8F",  -- 143
        12532 => X"88",  -- 136
        12533 => X"83",  -- 131
        12534 => X"80",  -- 128
        12535 => X"82",  -- 130
        12536 => X"83",  -- 131
        12537 => X"7A",  -- 122
        12538 => X"71",  -- 113
        12539 => X"6E",  -- 110
        12540 => X"6B",  -- 107
        12541 => X"67",  -- 103
        12542 => X"65",  -- 101
        12543 => X"68",  -- 104
        12544 => X"88",  -- 136
        12545 => X"7D",  -- 125
        12546 => X"69",  -- 105
        12547 => X"51",  -- 81
        12548 => X"3E",  -- 62
        12549 => X"32",  -- 50
        12550 => X"2A",  -- 42
        12551 => X"22",  -- 34
        12552 => X"13",  -- 19
        12553 => X"27",  -- 39
        12554 => X"41",  -- 65
        12555 => X"45",  -- 69
        12556 => X"50",  -- 80
        12557 => X"6A",  -- 106
        12558 => X"83",  -- 131
        12559 => X"82",  -- 130
        12560 => X"79",  -- 121
        12561 => X"8B",  -- 139
        12562 => X"7F",  -- 127
        12563 => X"7F",  -- 127
        12564 => X"7E",  -- 126
        12565 => X"73",  -- 115
        12566 => X"77",  -- 119
        12567 => X"6F",  -- 111
        12568 => X"66",  -- 102
        12569 => X"5D",  -- 93
        12570 => X"56",  -- 86
        12571 => X"37",  -- 55
        12572 => X"59",  -- 89
        12573 => X"57",  -- 87
        12574 => X"58",  -- 88
        12575 => X"3D",  -- 61
        12576 => X"20",  -- 32
        12577 => X"37",  -- 55
        12578 => X"42",  -- 66
        12579 => X"49",  -- 73
        12580 => X"45",  -- 69
        12581 => X"43",  -- 67
        12582 => X"56",  -- 86
        12583 => X"5D",  -- 93
        12584 => X"69",  -- 105
        12585 => X"66",  -- 102
        12586 => X"5C",  -- 92
        12587 => X"57",  -- 87
        12588 => X"61",  -- 97
        12589 => X"74",  -- 116
        12590 => X"7A",  -- 122
        12591 => X"77",  -- 119
        12592 => X"84",  -- 132
        12593 => X"91",  -- 145
        12594 => X"8D",  -- 141
        12595 => X"93",  -- 147
        12596 => X"8D",  -- 141
        12597 => X"89",  -- 137
        12598 => X"95",  -- 149
        12599 => X"7F",  -- 127
        12600 => X"81",  -- 129
        12601 => X"76",  -- 118
        12602 => X"74",  -- 116
        12603 => X"40",  -- 64
        12604 => X"26",  -- 38
        12605 => X"1D",  -- 29
        12606 => X"27",  -- 39
        12607 => X"28",  -- 40
        12608 => X"38",  -- 56
        12609 => X"48",  -- 72
        12610 => X"5E",  -- 94
        12611 => X"65",  -- 101
        12612 => X"71",  -- 113
        12613 => X"80",  -- 128
        12614 => X"77",  -- 119
        12615 => X"77",  -- 119
        12616 => X"55",  -- 85
        12617 => X"58",  -- 88
        12618 => X"67",  -- 103
        12619 => X"7B",  -- 123
        12620 => X"82",  -- 130
        12621 => X"7F",  -- 127
        12622 => X"7B",  -- 123
        12623 => X"7C",  -- 124
        12624 => X"7E",  -- 126
        12625 => X"85",  -- 133
        12626 => X"86",  -- 134
        12627 => X"7E",  -- 126
        12628 => X"7E",  -- 126
        12629 => X"86",  -- 134
        12630 => X"8B",  -- 139
        12631 => X"8B",  -- 139
        12632 => X"88",  -- 136
        12633 => X"88",  -- 136
        12634 => X"8A",  -- 138
        12635 => X"97",  -- 151
        12636 => X"A6",  -- 166
        12637 => X"AE",  -- 174
        12638 => X"A9",  -- 169
        12639 => X"A4",  -- 164
        12640 => X"A8",  -- 168
        12641 => X"B1",  -- 177
        12642 => X"B9",  -- 185
        12643 => X"BB",  -- 187
        12644 => X"B6",  -- 182
        12645 => X"B3",  -- 179
        12646 => X"B3",  -- 179
        12647 => X"B6",  -- 182
        12648 => X"B5",  -- 181
        12649 => X"AA",  -- 170
        12650 => X"A5",  -- 165
        12651 => X"A5",  -- 165
        12652 => X"9F",  -- 159
        12653 => X"88",  -- 136
        12654 => X"70",  -- 112
        12655 => X"62",  -- 98
        12656 => X"5E",  -- 94
        12657 => X"5D",  -- 93
        12658 => X"5B",  -- 91
        12659 => X"5A",  -- 90
        12660 => X"5D",  -- 93
        12661 => X"65",  -- 101
        12662 => X"6F",  -- 111
        12663 => X"78",  -- 120
        12664 => X"78",  -- 120
        12665 => X"73",  -- 115
        12666 => X"6F",  -- 111
        12667 => X"73",  -- 115
        12668 => X"79",  -- 121
        12669 => X"7E",  -- 126
        12670 => X"7F",  -- 127
        12671 => X"7D",  -- 125
        12672 => X"7C",  -- 124
        12673 => X"74",  -- 116
        12674 => X"77",  -- 119
        12675 => X"82",  -- 130
        12676 => X"83",  -- 131
        12677 => X"78",  -- 120
        12678 => X"73",  -- 115
        12679 => X"78",  -- 120
        12680 => X"71",  -- 113
        12681 => X"6C",  -- 108
        12682 => X"6C",  -- 108
        12683 => X"73",  -- 115
        12684 => X"7C",  -- 124
        12685 => X"80",  -- 128
        12686 => X"82",  -- 130
        12687 => X"84",  -- 132
        12688 => X"80",  -- 128
        12689 => X"80",  -- 128
        12690 => X"80",  -- 128
        12691 => X"7E",  -- 126
        12692 => X"7C",  -- 124
        12693 => X"80",  -- 128
        12694 => X"89",  -- 137
        12695 => X"90",  -- 144
        12696 => X"91",  -- 145
        12697 => X"95",  -- 149
        12698 => X"92",  -- 146
        12699 => X"8E",  -- 142
        12700 => X"92",  -- 146
        12701 => X"9B",  -- 155
        12702 => X"9B",  -- 155
        12703 => X"96",  -- 150
        12704 => X"9A",  -- 154
        12705 => X"9C",  -- 156
        12706 => X"9E",  -- 158
        12707 => X"9E",  -- 158
        12708 => X"9F",  -- 159
        12709 => X"A1",  -- 161
        12710 => X"9F",  -- 159
        12711 => X"9A",  -- 154
        12712 => X"98",  -- 152
        12713 => X"97",  -- 151
        12714 => X"94",  -- 148
        12715 => X"95",  -- 149
        12716 => X"96",  -- 150
        12717 => X"98",  -- 152
        12718 => X"99",  -- 153
        12719 => X"99",  -- 153
        12720 => X"88",  -- 136
        12721 => X"90",  -- 144
        12722 => X"8A",  -- 138
        12723 => X"79",  -- 121
        12724 => X"79",  -- 121
        12725 => X"8B",  -- 139
        12726 => X"97",  -- 151
        12727 => X"94",  -- 148
        12728 => X"92",  -- 146
        12729 => X"95",  -- 149
        12730 => X"9B",  -- 155
        12731 => X"A1",  -- 161
        12732 => X"A4",  -- 164
        12733 => X"A6",  -- 166
        12734 => X"A5",  -- 165
        12735 => X"A5",  -- 165
        12736 => X"A6",  -- 166
        12737 => X"A8",  -- 168
        12738 => X"AE",  -- 174
        12739 => X"B3",  -- 179
        12740 => X"B3",  -- 179
        12741 => X"AF",  -- 175
        12742 => X"A7",  -- 167
        12743 => X"A1",  -- 161
        12744 => X"9E",  -- 158
        12745 => X"9D",  -- 157
        12746 => X"9B",  -- 155
        12747 => X"98",  -- 152
        12748 => X"96",  -- 150
        12749 => X"97",  -- 151
        12750 => X"99",  -- 153
        12751 => X"9C",  -- 156
        12752 => X"92",  -- 146
        12753 => X"9A",  -- 154
        12754 => X"98",  -- 152
        12755 => X"7A",  -- 122
        12756 => X"51",  -- 81
        12757 => X"42",  -- 66
        12758 => X"40",  -- 64
        12759 => X"3B",  -- 59
        12760 => X"44",  -- 68
        12761 => X"61",  -- 97
        12762 => X"81",  -- 129
        12763 => X"90",  -- 144
        12764 => X"98",  -- 152
        12765 => X"9F",  -- 159
        12766 => X"A2",  -- 162
        12767 => X"9F",  -- 159
        12768 => X"96",  -- 150
        12769 => X"9C",  -- 156
        12770 => X"A3",  -- 163
        12771 => X"A7",  -- 167
        12772 => X"A9",  -- 169
        12773 => X"A2",  -- 162
        12774 => X"92",  -- 146
        12775 => X"83",  -- 131
        12776 => X"6E",  -- 110
        12777 => X"64",  -- 100
        12778 => X"5F",  -- 95
        12779 => X"6D",  -- 109
        12780 => X"89",  -- 137
        12781 => X"A1",  -- 161
        12782 => X"AF",  -- 175
        12783 => X"B1",  -- 177
        12784 => X"B4",  -- 180
        12785 => X"B2",  -- 178
        12786 => X"B0",  -- 176
        12787 => X"AE",  -- 174
        12788 => X"B1",  -- 177
        12789 => X"B6",  -- 182
        12790 => X"BD",  -- 189
        12791 => X"C1",  -- 193
        12792 => X"BF",  -- 191
        12793 => X"BB",  -- 187
        12794 => X"C1",  -- 193
        12795 => X"C4",  -- 196
        12796 => X"BD",  -- 189
        12797 => X"BF",  -- 191
        12798 => X"B8",  -- 184
        12799 => X"9E",  -- 158
        12800 => X"39",  -- 57
        12801 => X"3A",  -- 58
        12802 => X"3B",  -- 59
        12803 => X"3A",  -- 58
        12804 => X"3A",  -- 58
        12805 => X"3F",  -- 63
        12806 => X"45",  -- 69
        12807 => X"4A",  -- 74
        12808 => X"4A",  -- 74
        12809 => X"4E",  -- 78
        12810 => X"57",  -- 87
        12811 => X"5C",  -- 92
        12812 => X"60",  -- 96
        12813 => X"62",  -- 98
        12814 => X"66",  -- 102
        12815 => X"66",  -- 102
        12816 => X"6F",  -- 111
        12817 => X"6F",  -- 111
        12818 => X"6D",  -- 109
        12819 => X"6E",  -- 110
        12820 => X"76",  -- 118
        12821 => X"7E",  -- 126
        12822 => X"7B",  -- 123
        12823 => X"75",  -- 117
        12824 => X"72",  -- 114
        12825 => X"72",  -- 114
        12826 => X"6F",  -- 111
        12827 => X"67",  -- 103
        12828 => X"5E",  -- 94
        12829 => X"5A",  -- 90
        12830 => X"5B",  -- 91
        12831 => X"5E",  -- 94
        12832 => X"5E",  -- 94
        12833 => X"5E",  -- 94
        12834 => X"62",  -- 98
        12835 => X"66",  -- 102
        12836 => X"66",  -- 102
        12837 => X"64",  -- 100
        12838 => X"68",  -- 104
        12839 => X"6E",  -- 110
        12840 => X"76",  -- 118
        12841 => X"81",  -- 129
        12842 => X"88",  -- 136
        12843 => X"88",  -- 136
        12844 => X"8B",  -- 139
        12845 => X"94",  -- 148
        12846 => X"97",  -- 151
        12847 => X"95",  -- 149
        12848 => X"A5",  -- 165
        12849 => X"A2",  -- 162
        12850 => X"9D",  -- 157
        12851 => X"95",  -- 149
        12852 => X"8B",  -- 139
        12853 => X"85",  -- 133
        12854 => X"84",  -- 132
        12855 => X"82",  -- 130
        12856 => X"7E",  -- 126
        12857 => X"7D",  -- 125
        12858 => X"77",  -- 119
        12859 => X"7A",  -- 122
        12860 => X"71",  -- 113
        12861 => X"68",  -- 104
        12862 => X"6D",  -- 109
        12863 => X"61",  -- 97
        12864 => X"6C",  -- 108
        12865 => X"7A",  -- 122
        12866 => X"59",  -- 89
        12867 => X"47",  -- 71
        12868 => X"3B",  -- 59
        12869 => X"23",  -- 35
        12870 => X"24",  -- 36
        12871 => X"23",  -- 35
        12872 => X"2C",  -- 44
        12873 => X"45",  -- 69
        12874 => X"4B",  -- 75
        12875 => X"75",  -- 117
        12876 => X"7A",  -- 122
        12877 => X"81",  -- 129
        12878 => X"88",  -- 136
        12879 => X"88",  -- 136
        12880 => X"81",  -- 129
        12881 => X"82",  -- 130
        12882 => X"7B",  -- 123
        12883 => X"77",  -- 119
        12884 => X"77",  -- 119
        12885 => X"75",  -- 117
        12886 => X"65",  -- 101
        12887 => X"53",  -- 83
        12888 => X"3E",  -- 62
        12889 => X"36",  -- 54
        12890 => X"3E",  -- 62
        12891 => X"36",  -- 54
        12892 => X"30",  -- 48
        12893 => X"42",  -- 66
        12894 => X"3E",  -- 62
        12895 => X"2E",  -- 46
        12896 => X"22",  -- 34
        12897 => X"27",  -- 39
        12898 => X"29",  -- 41
        12899 => X"2B",  -- 43
        12900 => X"2D",  -- 45
        12901 => X"29",  -- 41
        12902 => X"2F",  -- 47
        12903 => X"42",  -- 66
        12904 => X"3F",  -- 63
        12905 => X"42",  -- 66
        12906 => X"35",  -- 53
        12907 => X"40",  -- 64
        12908 => X"48",  -- 72
        12909 => X"4C",  -- 76
        12910 => X"62",  -- 98
        12911 => X"61",  -- 97
        12912 => X"6F",  -- 111
        12913 => X"81",  -- 129
        12914 => X"92",  -- 146
        12915 => X"8B",  -- 139
        12916 => X"7F",  -- 127
        12917 => X"8A",  -- 138
        12918 => X"97",  -- 151
        12919 => X"93",  -- 147
        12920 => X"82",  -- 130
        12921 => X"94",  -- 148
        12922 => X"7C",  -- 124
        12923 => X"4E",  -- 78
        12924 => X"3F",  -- 63
        12925 => X"2B",  -- 43
        12926 => X"16",  -- 22
        12927 => X"31",  -- 49
        12928 => X"2E",  -- 46
        12929 => X"39",  -- 57
        12930 => X"41",  -- 65
        12931 => X"4B",  -- 75
        12932 => X"61",  -- 97
        12933 => X"5F",  -- 95
        12934 => X"86",  -- 134
        12935 => X"89",  -- 137
        12936 => X"6A",  -- 106
        12937 => X"68",  -- 104
        12938 => X"6C",  -- 108
        12939 => X"75",  -- 117
        12940 => X"7A",  -- 122
        12941 => X"76",  -- 118
        12942 => X"77",  -- 119
        12943 => X"7C",  -- 124
        12944 => X"84",  -- 132
        12945 => X"8A",  -- 138
        12946 => X"82",  -- 130
        12947 => X"83",  -- 131
        12948 => X"91",  -- 145
        12949 => X"90",  -- 144
        12950 => X"86",  -- 134
        12951 => X"8B",  -- 139
        12952 => X"93",  -- 147
        12953 => X"97",  -- 151
        12954 => X"A0",  -- 160
        12955 => X"A0",  -- 160
        12956 => X"9A",  -- 154
        12957 => X"9F",  -- 159
        12958 => X"A5",  -- 165
        12959 => X"A2",  -- 162
        12960 => X"A5",  -- 165
        12961 => X"A9",  -- 169
        12962 => X"B3",  -- 179
        12963 => X"BD",  -- 189
        12964 => X"BE",  -- 190
        12965 => X"B6",  -- 182
        12966 => X"B1",  -- 177
        12967 => X"B1",  -- 177
        12968 => X"B7",  -- 183
        12969 => X"B6",  -- 182
        12970 => X"A8",  -- 168
        12971 => X"95",  -- 149
        12972 => X"7F",  -- 127
        12973 => X"75",  -- 117
        12974 => X"77",  -- 119
        12975 => X"6E",  -- 110
        12976 => X"6E",  -- 110
        12977 => X"68",  -- 104
        12978 => X"61",  -- 97
        12979 => X"5E",  -- 94
        12980 => X"62",  -- 98
        12981 => X"65",  -- 101
        12982 => X"67",  -- 103
        12983 => X"67",  -- 103
        12984 => X"75",  -- 117
        12985 => X"76",  -- 118
        12986 => X"74",  -- 116
        12987 => X"70",  -- 112
        12988 => X"70",  -- 112
        12989 => X"74",  -- 116
        12990 => X"78",  -- 120
        12991 => X"77",  -- 119
        12992 => X"77",  -- 119
        12993 => X"7C",  -- 124
        12994 => X"7E",  -- 126
        12995 => X"7A",  -- 122
        12996 => X"77",  -- 119
        12997 => X"77",  -- 119
        12998 => X"74",  -- 116
        12999 => X"6F",  -- 111
        13000 => X"6D",  -- 109
        13001 => X"78",  -- 120
        13002 => X"81",  -- 129
        13003 => X"81",  -- 129
        13004 => X"80",  -- 128
        13005 => X"81",  -- 129
        13006 => X"81",  -- 129
        13007 => X"7F",  -- 127
        13008 => X"7E",  -- 126
        13009 => X"7B",  -- 123
        13010 => X"80",  -- 128
        13011 => X"85",  -- 133
        13012 => X"83",  -- 131
        13013 => X"7D",  -- 125
        13014 => X"83",  -- 131
        13015 => X"8E",  -- 142
        13016 => X"90",  -- 144
        13017 => X"98",  -- 152
        13018 => X"9B",  -- 155
        13019 => X"96",  -- 150
        13020 => X"91",  -- 145
        13021 => X"91",  -- 145
        13022 => X"93",  -- 147
        13023 => X"94",  -- 148
        13024 => X"9B",  -- 155
        13025 => X"9A",  -- 154
        13026 => X"9C",  -- 156
        13027 => X"A1",  -- 161
        13028 => X"A4",  -- 164
        13029 => X"A1",  -- 161
        13030 => X"9A",  -- 154
        13031 => X"92",  -- 146
        13032 => X"95",  -- 149
        13033 => X"93",  -- 147
        13034 => X"91",  -- 145
        13035 => X"92",  -- 146
        13036 => X"94",  -- 148
        13037 => X"94",  -- 148
        13038 => X"91",  -- 145
        13039 => X"8D",  -- 141
        13040 => X"87",  -- 135
        13041 => X"87",  -- 135
        13042 => X"86",  -- 134
        13043 => X"87",  -- 135
        13044 => X"90",  -- 144
        13045 => X"99",  -- 153
        13046 => X"9A",  -- 154
        13047 => X"97",  -- 151
        13048 => X"98",  -- 152
        13049 => X"97",  -- 151
        13050 => X"97",  -- 151
        13051 => X"99",  -- 153
        13052 => X"9D",  -- 157
        13053 => X"A1",  -- 161
        13054 => X"A6",  -- 166
        13055 => X"AA",  -- 170
        13056 => X"A6",  -- 166
        13057 => X"A5",  -- 165
        13058 => X"AA",  -- 170
        13059 => X"B3",  -- 179
        13060 => X"B6",  -- 182
        13061 => X"B0",  -- 176
        13062 => X"A9",  -- 169
        13063 => X"A7",  -- 167
        13064 => X"9F",  -- 159
        13065 => X"A0",  -- 160
        13066 => X"9E",  -- 158
        13067 => X"9A",  -- 154
        13068 => X"97",  -- 151
        13069 => X"97",  -- 151
        13070 => X"98",  -- 152
        13071 => X"9A",  -- 154
        13072 => X"95",  -- 149
        13073 => X"97",  -- 151
        13074 => X"94",  -- 148
        13075 => X"83",  -- 131
        13076 => X"66",  -- 102
        13077 => X"49",  -- 73
        13078 => X"3E",  -- 62
        13079 => X"41",  -- 65
        13080 => X"4F",  -- 79
        13081 => X"5E",  -- 94
        13082 => X"78",  -- 120
        13083 => X"92",  -- 146
        13084 => X"9D",  -- 157
        13085 => X"9F",  -- 159
        13086 => X"9F",  -- 159
        13087 => X"A2",  -- 162
        13088 => X"A1",  -- 161
        13089 => X"A1",  -- 161
        13090 => X"A6",  -- 166
        13091 => X"A4",  -- 164
        13092 => X"A1",  -- 161
        13093 => X"A1",  -- 161
        13094 => X"99",  -- 153
        13095 => X"86",  -- 134
        13096 => X"71",  -- 113
        13097 => X"5E",  -- 94
        13098 => X"5E",  -- 94
        13099 => X"77",  -- 119
        13100 => X"93",  -- 147
        13101 => X"A8",  -- 168
        13102 => X"B2",  -- 178
        13103 => X"AD",  -- 173
        13104 => X"AD",  -- 173
        13105 => X"B1",  -- 177
        13106 => X"B6",  -- 182
        13107 => X"B2",  -- 178
        13108 => X"AD",  -- 173
        13109 => X"AF",  -- 175
        13110 => X"BB",  -- 187
        13111 => X"C5",  -- 197
        13112 => X"BC",  -- 188
        13113 => X"C2",  -- 194
        13114 => X"C3",  -- 195
        13115 => X"B8",  -- 184
        13116 => X"C1",  -- 193
        13117 => X"C7",  -- 199
        13118 => X"AB",  -- 171
        13119 => X"9A",  -- 154
        13120 => X"3C",  -- 60
        13121 => X"3F",  -- 63
        13122 => X"43",  -- 67
        13123 => X"45",  -- 69
        13124 => X"49",  -- 73
        13125 => X"4D",  -- 77
        13126 => X"52",  -- 82
        13127 => X"58",  -- 88
        13128 => X"61",  -- 97
        13129 => X"67",  -- 103
        13130 => X"6E",  -- 110
        13131 => X"76",  -- 118
        13132 => X"7B",  -- 123
        13133 => X"7B",  -- 123
        13134 => X"7A",  -- 122
        13135 => X"7A",  -- 122
        13136 => X"77",  -- 119
        13137 => X"78",  -- 120
        13138 => X"75",  -- 117
        13139 => X"71",  -- 113
        13140 => X"72",  -- 114
        13141 => X"76",  -- 118
        13142 => X"75",  -- 117
        13143 => X"70",  -- 112
        13144 => X"69",  -- 105
        13145 => X"6B",  -- 107
        13146 => X"69",  -- 105
        13147 => X"64",  -- 100
        13148 => X"5E",  -- 94
        13149 => X"58",  -- 88
        13150 => X"59",  -- 89
        13151 => X"5A",  -- 90
        13152 => X"5E",  -- 94
        13153 => X"5E",  -- 94
        13154 => X"61",  -- 97
        13155 => X"68",  -- 104
        13156 => X"70",  -- 112
        13157 => X"75",  -- 117
        13158 => X"77",  -- 119
        13159 => X"76",  -- 118
        13160 => X"86",  -- 134
        13161 => X"7E",  -- 126
        13162 => X"83",  -- 131
        13163 => X"94",  -- 148
        13164 => X"97",  -- 151
        13165 => X"8E",  -- 142
        13166 => X"91",  -- 145
        13167 => X"9E",  -- 158
        13168 => X"97",  -- 151
        13169 => X"98",  -- 152
        13170 => X"9A",  -- 154
        13171 => X"98",  -- 152
        13172 => X"93",  -- 147
        13173 => X"8B",  -- 139
        13174 => X"83",  -- 131
        13175 => X"7F",  -- 127
        13176 => X"7A",  -- 122
        13177 => X"76",  -- 118
        13178 => X"6E",  -- 110
        13179 => X"77",  -- 119
        13180 => X"78",  -- 120
        13181 => X"75",  -- 117
        13182 => X"75",  -- 117
        13183 => X"64",  -- 100
        13184 => X"53",  -- 83
        13185 => X"55",  -- 85
        13186 => X"3A",  -- 58
        13187 => X"2A",  -- 42
        13188 => X"27",  -- 39
        13189 => X"21",  -- 33
        13190 => X"29",  -- 41
        13191 => X"35",  -- 53
        13192 => X"5B",  -- 91
        13193 => X"6C",  -- 108
        13194 => X"72",  -- 114
        13195 => X"7D",  -- 125
        13196 => X"81",  -- 129
        13197 => X"78",  -- 120
        13198 => X"89",  -- 137
        13199 => X"86",  -- 134
        13200 => X"7D",  -- 125
        13201 => X"7F",  -- 127
        13202 => X"7F",  -- 127
        13203 => X"79",  -- 121
        13204 => X"6E",  -- 110
        13205 => X"5E",  -- 94
        13206 => X"46",  -- 70
        13207 => X"34",  -- 52
        13208 => X"2C",  -- 44
        13209 => X"1D",  -- 29
        13210 => X"1E",  -- 30
        13211 => X"1C",  -- 28
        13212 => X"26",  -- 38
        13213 => X"37",  -- 55
        13214 => X"29",  -- 41
        13215 => X"18",  -- 24
        13216 => X"1E",  -- 30
        13217 => X"22",  -- 34
        13218 => X"1F",  -- 31
        13219 => X"1F",  -- 31
        13220 => X"25",  -- 37
        13221 => X"24",  -- 36
        13222 => X"23",  -- 35
        13223 => X"2E",  -- 46
        13224 => X"27",  -- 39
        13225 => X"2B",  -- 43
        13226 => X"28",  -- 40
        13227 => X"38",  -- 56
        13228 => X"39",  -- 57
        13229 => X"2C",  -- 44
        13230 => X"37",  -- 55
        13231 => X"38",  -- 56
        13232 => X"4E",  -- 78
        13233 => X"5E",  -- 94
        13234 => X"74",  -- 116
        13235 => X"78",  -- 120
        13236 => X"77",  -- 119
        13237 => X"84",  -- 132
        13238 => X"90",  -- 144
        13239 => X"8C",  -- 140
        13240 => X"92",  -- 146
        13241 => X"8B",  -- 139
        13242 => X"80",  -- 128
        13243 => X"75",  -- 117
        13244 => X"5C",  -- 92
        13245 => X"36",  -- 54
        13246 => X"23",  -- 35
        13247 => X"1F",  -- 31
        13248 => X"24",  -- 36
        13249 => X"2D",  -- 45
        13250 => X"38",  -- 56
        13251 => X"42",  -- 66
        13252 => X"4C",  -- 76
        13253 => X"40",  -- 64
        13254 => X"67",  -- 103
        13255 => X"77",  -- 119
        13256 => X"74",  -- 116
        13257 => X"73",  -- 115
        13258 => X"77",  -- 119
        13259 => X"7C",  -- 124
        13260 => X"7F",  -- 127
        13261 => X"7C",  -- 124
        13262 => X"7A",  -- 122
        13263 => X"7B",  -- 123
        13264 => X"7F",  -- 127
        13265 => X"81",  -- 129
        13266 => X"80",  -- 128
        13267 => X"81",  -- 129
        13268 => X"8A",  -- 138
        13269 => X"8C",  -- 140
        13270 => X"8B",  -- 139
        13271 => X"90",  -- 144
        13272 => X"91",  -- 145
        13273 => X"95",  -- 149
        13274 => X"9A",  -- 154
        13275 => X"9D",  -- 157
        13276 => X"9C",  -- 156
        13277 => X"99",  -- 153
        13278 => X"97",  -- 151
        13279 => X"97",  -- 151
        13280 => X"9C",  -- 156
        13281 => X"8E",  -- 142
        13282 => X"92",  -- 146
        13283 => X"AB",  -- 171
        13284 => X"BC",  -- 188
        13285 => X"BB",  -- 187
        13286 => X"BC",  -- 188
        13287 => X"C8",  -- 200
        13288 => X"BC",  -- 188
        13289 => X"B3",  -- 179
        13290 => X"BA",  -- 186
        13291 => X"AE",  -- 174
        13292 => X"7D",  -- 125
        13293 => X"6D",  -- 109
        13294 => X"78",  -- 120
        13295 => X"68",  -- 104
        13296 => X"66",  -- 102
        13297 => X"61",  -- 97
        13298 => X"5C",  -- 92
        13299 => X"5D",  -- 93
        13300 => X"61",  -- 97
        13301 => X"66",  -- 102
        13302 => X"66",  -- 102
        13303 => X"65",  -- 101
        13304 => X"65",  -- 101
        13305 => X"65",  -- 101
        13306 => X"62",  -- 98
        13307 => X"5F",  -- 95
        13308 => X"62",  -- 98
        13309 => X"68",  -- 104
        13310 => X"6C",  -- 108
        13311 => X"6C",  -- 108
        13312 => X"71",  -- 113
        13313 => X"72",  -- 114
        13314 => X"72",  -- 114
        13315 => X"70",  -- 112
        13316 => X"73",  -- 115
        13317 => X"76",  -- 118
        13318 => X"74",  -- 116
        13319 => X"6E",  -- 110
        13320 => X"7A",  -- 122
        13321 => X"7D",  -- 125
        13322 => X"7C",  -- 124
        13323 => X"79",  -- 121
        13324 => X"7A",  -- 122
        13325 => X"7E",  -- 126
        13326 => X"80",  -- 128
        13327 => X"7F",  -- 127
        13328 => X"81",  -- 129
        13329 => X"80",  -- 128
        13330 => X"85",  -- 133
        13331 => X"8B",  -- 139
        13332 => X"86",  -- 134
        13333 => X"7C",  -- 124
        13334 => X"7C",  -- 124
        13335 => X"82",  -- 130
        13336 => X"92",  -- 146
        13337 => X"98",  -- 152
        13338 => X"9A",  -- 154
        13339 => X"97",  -- 151
        13340 => X"95",  -- 149
        13341 => X"96",  -- 150
        13342 => X"97",  -- 151
        13343 => X"97",  -- 151
        13344 => X"9C",  -- 156
        13345 => X"9C",  -- 156
        13346 => X"9D",  -- 157
        13347 => X"9F",  -- 159
        13348 => X"9E",  -- 158
        13349 => X"9A",  -- 154
        13350 => X"94",  -- 148
        13351 => X"8F",  -- 143
        13352 => X"92",  -- 146
        13353 => X"91",  -- 145
        13354 => X"8F",  -- 143
        13355 => X"90",  -- 144
        13356 => X"91",  -- 145
        13357 => X"90",  -- 144
        13358 => X"8F",  -- 143
        13359 => X"8D",  -- 141
        13360 => X"8E",  -- 142
        13361 => X"87",  -- 135
        13362 => X"88",  -- 136
        13363 => X"8F",  -- 143
        13364 => X"90",  -- 144
        13365 => X"8A",  -- 138
        13366 => X"8E",  -- 142
        13367 => X"9B",  -- 155
        13368 => X"96",  -- 150
        13369 => X"97",  -- 151
        13370 => X"99",  -- 153
        13371 => X"9D",  -- 157
        13372 => X"A0",  -- 160
        13373 => X"A3",  -- 163
        13374 => X"A7",  -- 167
        13375 => X"AB",  -- 171
        13376 => X"A0",  -- 160
        13377 => X"A0",  -- 160
        13378 => X"A5",  -- 165
        13379 => X"AE",  -- 174
        13380 => X"B2",  -- 178
        13381 => X"AF",  -- 175
        13382 => X"AA",  -- 170
        13383 => X"A9",  -- 169
        13384 => X"9D",  -- 157
        13385 => X"9C",  -- 156
        13386 => X"99",  -- 153
        13387 => X"95",  -- 149
        13388 => X"94",  -- 148
        13389 => X"94",  -- 148
        13390 => X"96",  -- 150
        13391 => X"97",  -- 151
        13392 => X"94",  -- 148
        13393 => X"99",  -- 153
        13394 => X"97",  -- 151
        13395 => X"80",  -- 128
        13396 => X"5D",  -- 93
        13397 => X"45",  -- 69
        13398 => X"45",  -- 69
        13399 => X"51",  -- 81
        13400 => X"56",  -- 86
        13401 => X"61",  -- 97
        13402 => X"73",  -- 115
        13403 => X"86",  -- 134
        13404 => X"8F",  -- 143
        13405 => X"92",  -- 146
        13406 => X"96",  -- 150
        13407 => X"9C",  -- 156
        13408 => X"9E",  -- 158
        13409 => X"9E",  -- 158
        13410 => X"A1",  -- 161
        13411 => X"A0",  -- 160
        13412 => X"9D",  -- 157
        13413 => X"A0",  -- 160
        13414 => X"99",  -- 153
        13415 => X"88",  -- 136
        13416 => X"7C",  -- 124
        13417 => X"68",  -- 104
        13418 => X"69",  -- 105
        13419 => X"81",  -- 129
        13420 => X"9B",  -- 155
        13421 => X"AC",  -- 172
        13422 => X"B1",  -- 177
        13423 => X"A8",  -- 168
        13424 => X"A9",  -- 169
        13425 => X"AE",  -- 174
        13426 => X"B1",  -- 177
        13427 => X"B1",  -- 177
        13428 => X"AF",  -- 175
        13429 => X"B2",  -- 178
        13430 => X"BC",  -- 188
        13431 => X"C4",  -- 196
        13432 => X"C6",  -- 198
        13433 => X"C6",  -- 198
        13434 => X"C4",  -- 196
        13435 => X"BA",  -- 186
        13436 => X"C0",  -- 192
        13437 => X"BD",  -- 189
        13438 => X"9D",  -- 157
        13439 => X"8C",  -- 140
        13440 => X"4F",  -- 79
        13441 => X"54",  -- 84
        13442 => X"59",  -- 89
        13443 => X"5F",  -- 95
        13444 => X"61",  -- 97
        13445 => X"66",  -- 102
        13446 => X"68",  -- 104
        13447 => X"6B",  -- 107
        13448 => X"72",  -- 114
        13449 => X"74",  -- 116
        13450 => X"7A",  -- 122
        13451 => X"82",  -- 130
        13452 => X"88",  -- 136
        13453 => X"8A",  -- 138
        13454 => X"86",  -- 134
        13455 => X"82",  -- 130
        13456 => X"7B",  -- 123
        13457 => X"7B",  -- 123
        13458 => X"76",  -- 118
        13459 => X"6F",  -- 111
        13460 => X"6C",  -- 108
        13461 => X"6D",  -- 109
        13462 => X"70",  -- 112
        13463 => X"71",  -- 113
        13464 => X"65",  -- 101
        13465 => X"69",  -- 105
        13466 => X"6C",  -- 108
        13467 => X"6B",  -- 107
        13468 => X"67",  -- 103
        13469 => X"63",  -- 99
        13470 => X"65",  -- 101
        13471 => X"66",  -- 102
        13472 => X"6B",  -- 107
        13473 => X"74",  -- 116
        13474 => X"7A",  -- 122
        13475 => X"75",  -- 117
        13476 => X"70",  -- 112
        13477 => X"74",  -- 116
        13478 => X"76",  -- 118
        13479 => X"73",  -- 115
        13480 => X"7F",  -- 127
        13481 => X"86",  -- 134
        13482 => X"8B",  -- 139
        13483 => X"90",  -- 144
        13484 => X"97",  -- 151
        13485 => X"9C",  -- 156
        13486 => X"99",  -- 153
        13487 => X"93",  -- 147
        13488 => X"94",  -- 148
        13489 => X"93",  -- 147
        13490 => X"93",  -- 147
        13491 => X"94",  -- 148
        13492 => X"92",  -- 146
        13493 => X"8D",  -- 141
        13494 => X"86",  -- 134
        13495 => X"81",  -- 129
        13496 => X"7E",  -- 126
        13497 => X"7E",  -- 126
        13498 => X"71",  -- 113
        13499 => X"6E",  -- 110
        13500 => X"66",  -- 102
        13501 => X"54",  -- 84
        13502 => X"4D",  -- 77
        13503 => X"3C",  -- 60
        13504 => X"39",  -- 57
        13505 => X"33",  -- 51
        13506 => X"2F",  -- 47
        13507 => X"2B",  -- 43
        13508 => X"32",  -- 50
        13509 => X"3C",  -- 60
        13510 => X"43",  -- 67
        13511 => X"5B",  -- 91
        13512 => X"78",  -- 120
        13513 => X"7B",  -- 123
        13514 => X"81",  -- 129
        13515 => X"7A",  -- 122
        13516 => X"88",  -- 136
        13517 => X"7B",  -- 123
        13518 => X"84",  -- 132
        13519 => X"73",  -- 115
        13520 => X"66",  -- 102
        13521 => X"60",  -- 96
        13522 => X"5A",  -- 90
        13523 => X"52",  -- 82
        13524 => X"44",  -- 68
        13525 => X"37",  -- 55
        13526 => X"2E",  -- 46
        13527 => X"2D",  -- 45
        13528 => X"25",  -- 37
        13529 => X"17",  -- 23
        13530 => X"12",  -- 18
        13531 => X"11",  -- 17
        13532 => X"26",  -- 38
        13533 => X"34",  -- 52
        13534 => X"27",  -- 39
        13535 => X"27",  -- 39
        13536 => X"16",  -- 22
        13537 => X"1C",  -- 28
        13538 => X"18",  -- 24
        13539 => X"18",  -- 24
        13540 => X"23",  -- 35
        13541 => X"26",  -- 38
        13542 => X"20",  -- 32
        13543 => X"1D",  -- 29
        13544 => X"18",  -- 24
        13545 => X"24",  -- 36
        13546 => X"26",  -- 38
        13547 => X"30",  -- 48
        13548 => X"2B",  -- 43
        13549 => X"1F",  -- 31
        13550 => X"23",  -- 35
        13551 => X"23",  -- 35
        13552 => X"33",  -- 51
        13553 => X"35",  -- 53
        13554 => X"40",  -- 64
        13555 => X"46",  -- 70
        13556 => X"4E",  -- 78
        13557 => X"68",  -- 104
        13558 => X"82",  -- 130
        13559 => X"8C",  -- 140
        13560 => X"8D",  -- 141
        13561 => X"83",  -- 131
        13562 => X"84",  -- 132
        13563 => X"8D",  -- 141
        13564 => X"6D",  -- 109
        13565 => X"52",  -- 82
        13566 => X"49",  -- 73
        13567 => X"1B",  -- 27
        13568 => X"25",  -- 37
        13569 => X"33",  -- 51
        13570 => X"45",  -- 69
        13571 => X"51",  -- 81
        13572 => X"4E",  -- 78
        13573 => X"3B",  -- 59
        13574 => X"57",  -- 87
        13575 => X"6F",  -- 111
        13576 => X"72",  -- 114
        13577 => X"73",  -- 115
        13578 => X"74",  -- 116
        13579 => X"77",  -- 119
        13580 => X"7B",  -- 123
        13581 => X"7F",  -- 127
        13582 => X"7F",  -- 127
        13583 => X"7A",  -- 122
        13584 => X"86",  -- 134
        13585 => X"7F",  -- 127
        13586 => X"82",  -- 130
        13587 => X"88",  -- 136
        13588 => X"8B",  -- 139
        13589 => X"87",  -- 135
        13590 => X"79",  -- 121
        13591 => X"66",  -- 102
        13592 => X"7A",  -- 122
        13593 => X"7E",  -- 126
        13594 => X"7D",  -- 125
        13595 => X"82",  -- 130
        13596 => X"87",  -- 135
        13597 => X"6E",  -- 110
        13598 => X"4C",  -- 76
        13599 => X"45",  -- 69
        13600 => X"38",  -- 56
        13601 => X"28",  -- 40
        13602 => X"31",  -- 49
        13603 => X"5B",  -- 91
        13604 => X"7E",  -- 126
        13605 => X"88",  -- 136
        13606 => X"9D",  -- 157
        13607 => X"BB",  -- 187
        13608 => X"BE",  -- 190
        13609 => X"C4",  -- 196
        13610 => X"B8",  -- 184
        13611 => X"AB",  -- 171
        13612 => X"AB",  -- 171
        13613 => X"99",  -- 153
        13614 => X"7E",  -- 126
        13615 => X"73",  -- 115
        13616 => X"6C",  -- 108
        13617 => X"67",  -- 103
        13618 => X"64",  -- 100
        13619 => X"65",  -- 101
        13620 => X"6B",  -- 107
        13621 => X"6F",  -- 111
        13622 => X"6F",  -- 111
        13623 => X"6C",  -- 108
        13624 => X"62",  -- 98
        13625 => X"64",  -- 100
        13626 => X"64",  -- 100
        13627 => X"65",  -- 101
        13628 => X"69",  -- 105
        13629 => X"6F",  -- 111
        13630 => X"70",  -- 112
        13631 => X"6D",  -- 109
        13632 => X"6C",  -- 108
        13633 => X"6A",  -- 106
        13634 => X"6A",  -- 106
        13635 => X"6C",  -- 108
        13636 => X"74",  -- 116
        13637 => X"7A",  -- 122
        13638 => X"7A",  -- 122
        13639 => X"75",  -- 117
        13640 => X"7C",  -- 124
        13641 => X"7B",  -- 123
        13642 => X"76",  -- 118
        13643 => X"74",  -- 116
        13644 => X"77",  -- 119
        13645 => X"7C",  -- 124
        13646 => X"7D",  -- 125
        13647 => X"7B",  -- 123
        13648 => X"7D",  -- 125
        13649 => X"7E",  -- 126
        13650 => X"84",  -- 132
        13651 => X"8A",  -- 138
        13652 => X"85",  -- 133
        13653 => X"78",  -- 120
        13654 => X"72",  -- 114
        13655 => X"72",  -- 114
        13656 => X"87",  -- 135
        13657 => X"8C",  -- 140
        13658 => X"8F",  -- 143
        13659 => X"8F",  -- 143
        13660 => X"90",  -- 144
        13661 => X"92",  -- 146
        13662 => X"93",  -- 147
        13663 => X"93",  -- 147
        13664 => X"9D",  -- 157
        13665 => X"9F",  -- 159
        13666 => X"9F",  -- 159
        13667 => X"9E",  -- 158
        13668 => X"99",  -- 153
        13669 => X"95",  -- 149
        13670 => X"92",  -- 146
        13671 => X"90",  -- 144
        13672 => X"90",  -- 144
        13673 => X"8F",  -- 143
        13674 => X"8D",  -- 141
        13675 => X"8B",  -- 139
        13676 => X"89",  -- 137
        13677 => X"87",  -- 135
        13678 => X"87",  -- 135
        13679 => X"85",  -- 133
        13680 => X"8B",  -- 139
        13681 => X"8B",  -- 139
        13682 => X"90",  -- 144
        13683 => X"8F",  -- 143
        13684 => X"85",  -- 133
        13685 => X"7F",  -- 127
        13686 => X"88",  -- 136
        13687 => X"99",  -- 153
        13688 => X"93",  -- 147
        13689 => X"97",  -- 151
        13690 => X"9A",  -- 154
        13691 => X"9D",  -- 157
        13692 => X"A0",  -- 160
        13693 => X"A3",  -- 163
        13694 => X"A5",  -- 165
        13695 => X"A8",  -- 168
        13696 => X"9E",  -- 158
        13697 => X"9E",  -- 158
        13698 => X"A3",  -- 163
        13699 => X"AA",  -- 170
        13700 => X"AE",  -- 174
        13701 => X"AC",  -- 172
        13702 => X"AA",  -- 170
        13703 => X"A9",  -- 169
        13704 => X"9F",  -- 159
        13705 => X"99",  -- 153
        13706 => X"95",  -- 149
        13707 => X"92",  -- 146
        13708 => X"95",  -- 149
        13709 => X"96",  -- 150
        13710 => X"97",  -- 151
        13711 => X"98",  -- 152
        13712 => X"9A",  -- 154
        13713 => X"9C",  -- 156
        13714 => X"96",  -- 150
        13715 => X"82",  -- 130
        13716 => X"65",  -- 101
        13717 => X"4F",  -- 79
        13718 => X"4D",  -- 77
        13719 => X"57",  -- 87
        13720 => X"45",  -- 69
        13721 => X"4F",  -- 79
        13722 => X"62",  -- 98
        13723 => X"76",  -- 118
        13724 => X"84",  -- 132
        13725 => X"8B",  -- 139
        13726 => X"92",  -- 146
        13727 => X"98",  -- 152
        13728 => X"9C",  -- 156
        13729 => X"9B",  -- 155
        13730 => X"9D",  -- 157
        13731 => X"9C",  -- 156
        13732 => X"9A",  -- 154
        13733 => X"9E",  -- 158
        13734 => X"9A",  -- 154
        13735 => X"8A",  -- 138
        13736 => X"7A",  -- 122
        13737 => X"62",  -- 98
        13738 => X"5E",  -- 94
        13739 => X"76",  -- 118
        13740 => X"91",  -- 145
        13741 => X"A2",  -- 162
        13742 => X"A6",  -- 166
        13743 => X"9E",  -- 158
        13744 => X"A6",  -- 166
        13745 => X"A9",  -- 169
        13746 => X"AC",  -- 172
        13747 => X"AE",  -- 174
        13748 => X"B1",  -- 177
        13749 => X"B6",  -- 182
        13750 => X"BE",  -- 190
        13751 => X"C4",  -- 196
        13752 => X"C5",  -- 197
        13753 => X"C1",  -- 193
        13754 => X"C1",  -- 193
        13755 => X"BE",  -- 190
        13756 => X"C4",  -- 196
        13757 => X"B8",  -- 184
        13758 => X"97",  -- 151
        13759 => X"8D",  -- 141
        13760 => X"66",  -- 102
        13761 => X"6A",  -- 106
        13762 => X"6F",  -- 111
        13763 => X"74",  -- 116
        13764 => X"75",  -- 117
        13765 => X"74",  -- 116
        13766 => X"72",  -- 114
        13767 => X"71",  -- 113
        13768 => X"6F",  -- 111
        13769 => X"70",  -- 112
        13770 => X"73",  -- 115
        13771 => X"7B",  -- 123
        13772 => X"82",  -- 130
        13773 => X"85",  -- 133
        13774 => X"80",  -- 128
        13775 => X"7C",  -- 124
        13776 => X"7B",  -- 123
        13777 => X"78",  -- 120
        13778 => X"73",  -- 115
        13779 => X"6E",  -- 110
        13780 => X"6E",  -- 110
        13781 => X"71",  -- 113
        13782 => X"74",  -- 116
        13783 => X"75",  -- 117
        13784 => X"70",  -- 112
        13785 => X"73",  -- 115
        13786 => X"73",  -- 115
        13787 => X"6E",  -- 110
        13788 => X"67",  -- 103
        13789 => X"62",  -- 98
        13790 => X"62",  -- 98
        13791 => X"63",  -- 99
        13792 => X"6D",  -- 109
        13793 => X"7D",  -- 125
        13794 => X"88",  -- 136
        13795 => X"85",  -- 133
        13796 => X"84",  -- 132
        13797 => X"87",  -- 135
        13798 => X"84",  -- 132
        13799 => X"7A",  -- 122
        13800 => X"75",  -- 117
        13801 => X"7D",  -- 125
        13802 => X"7E",  -- 126
        13803 => X"7C",  -- 124
        13804 => X"87",  -- 135
        13805 => X"97",  -- 151
        13806 => X"90",  -- 144
        13807 => X"7E",  -- 126
        13808 => X"83",  -- 131
        13809 => X"85",  -- 133
        13810 => X"88",  -- 136
        13811 => X"8C",  -- 140
        13812 => X"8E",  -- 142
        13813 => X"8C",  -- 140
        13814 => X"87",  -- 135
        13815 => X"83",  -- 131
        13816 => X"7A",  -- 122
        13817 => X"88",  -- 136
        13818 => X"7E",  -- 126
        13819 => X"6E",  -- 110
        13820 => X"56",  -- 86
        13821 => X"3E",  -- 62
        13822 => X"3C",  -- 60
        13823 => X"3B",  -- 59
        13824 => X"37",  -- 55
        13825 => X"34",  -- 52
        13826 => X"48",  -- 72
        13827 => X"4E",  -- 78
        13828 => X"56",  -- 86
        13829 => X"60",  -- 96
        13830 => X"5C",  -- 92
        13831 => X"76",  -- 118
        13832 => X"74",  -- 116
        13833 => X"7A",  -- 122
        13834 => X"7E",  -- 126
        13835 => X"74",  -- 116
        13836 => X"79",  -- 121
        13837 => X"6C",  -- 108
        13838 => X"68",  -- 104
        13839 => X"54",  -- 84
        13840 => X"3B",  -- 59
        13841 => X"2D",  -- 45
        13842 => X"22",  -- 34
        13843 => X"1C",  -- 28
        13844 => X"16",  -- 22
        13845 => X"15",  -- 21
        13846 => X"1C",  -- 28
        13847 => X"29",  -- 41
        13848 => X"19",  -- 25
        13849 => X"15",  -- 21
        13850 => X"10",  -- 16
        13851 => X"0D",  -- 13
        13852 => X"1C",  -- 28
        13853 => X"27",  -- 39
        13854 => X"2D",  -- 45
        13855 => X"4A",  -- 74
        13856 => X"22",  -- 34
        13857 => X"29",  -- 41
        13858 => X"24",  -- 36
        13859 => X"1E",  -- 30
        13860 => X"24",  -- 36
        13861 => X"26",  -- 38
        13862 => X"1D",  -- 29
        13863 => X"16",  -- 22
        13864 => X"16",  -- 22
        13865 => X"21",  -- 33
        13866 => X"22",  -- 34
        13867 => X"1A",  -- 26
        13868 => X"16",  -- 22
        13869 => X"1B",  -- 27
        13870 => X"20",  -- 32
        13871 => X"1D",  -- 29
        13872 => X"27",  -- 39
        13873 => X"1F",  -- 31
        13874 => X"1D",  -- 29
        13875 => X"20",  -- 32
        13876 => X"28",  -- 40
        13877 => X"42",  -- 66
        13878 => X"65",  -- 101
        13879 => X"76",  -- 118
        13880 => X"70",  -- 112
        13881 => X"8A",  -- 138
        13882 => X"8A",  -- 138
        13883 => X"88",  -- 136
        13884 => X"71",  -- 113
        13885 => X"71",  -- 113
        13886 => X"71",  -- 113
        13887 => X"28",  -- 40
        13888 => X"22",  -- 34
        13889 => X"30",  -- 48
        13890 => X"44",  -- 68
        13891 => X"4E",  -- 78
        13892 => X"4B",  -- 75
        13893 => X"44",  -- 68
        13894 => X"56",  -- 86
        13895 => X"69",  -- 105
        13896 => X"68",  -- 104
        13897 => X"6E",  -- 110
        13898 => X"6F",  -- 111
        13899 => X"70",  -- 112
        13900 => X"75",  -- 117
        13901 => X"7C",  -- 124
        13902 => X"7B",  -- 123
        13903 => X"73",  -- 115
        13904 => X"6D",  -- 109
        13905 => X"65",  -- 101
        13906 => X"64",  -- 100
        13907 => X"57",  -- 87
        13908 => X"3D",  -- 61
        13909 => X"3D",  -- 61
        13910 => X"4F",  -- 79
        13911 => X"54",  -- 84
        13912 => X"67",  -- 103
        13913 => X"64",  -- 100
        13914 => X"48",  -- 72
        13915 => X"2B",  -- 43
        13916 => X"22",  -- 34
        13917 => X"17",  -- 23
        13918 => X"27",  -- 39
        13919 => X"53",  -- 83
        13920 => X"4D",  -- 77
        13921 => X"45",  -- 69
        13922 => X"42",  -- 66
        13923 => X"33",  -- 51
        13924 => X"14",  -- 20
        13925 => X"08",  -- 8
        13926 => X"2C",  -- 44
        13927 => X"6A",  -- 106
        13928 => X"B1",  -- 177
        13929 => X"C0",  -- 192
        13930 => X"BC",  -- 188
        13931 => X"A9",  -- 169
        13932 => X"A6",  -- 166
        13933 => X"97",  -- 151
        13934 => X"78",  -- 120
        13935 => X"73",  -- 115
        13936 => X"6D",  -- 109
        13937 => X"68",  -- 104
        13938 => X"63",  -- 99
        13939 => X"62",  -- 98
        13940 => X"66",  -- 102
        13941 => X"69",  -- 105
        13942 => X"68",  -- 104
        13943 => X"66",  -- 102
        13944 => X"68",  -- 104
        13945 => X"6B",  -- 107
        13946 => X"71",  -- 113
        13947 => X"75",  -- 117
        13948 => X"7B",  -- 123
        13949 => X"7D",  -- 125
        13950 => X"79",  -- 121
        13951 => X"71",  -- 113
        13952 => X"6B",  -- 107
        13953 => X"69",  -- 105
        13954 => X"6B",  -- 107
        13955 => X"6F",  -- 111
        13956 => X"75",  -- 117
        13957 => X"7A",  -- 122
        13958 => X"7B",  -- 123
        13959 => X"79",  -- 121
        13960 => X"74",  -- 116
        13961 => X"76",  -- 118
        13962 => X"78",  -- 120
        13963 => X"7A",  -- 122
        13964 => X"7D",  -- 125
        13965 => X"7E",  -- 126
        13966 => X"7C",  -- 124
        13967 => X"7A",  -- 122
        13968 => X"79",  -- 121
        13969 => X"7B",  -- 123
        13970 => X"81",  -- 129
        13971 => X"87",  -- 135
        13972 => X"84",  -- 132
        13973 => X"79",  -- 121
        13974 => X"72",  -- 114
        13975 => X"70",  -- 112
        13976 => X"79",  -- 121
        13977 => X"7F",  -- 127
        13978 => X"85",  -- 133
        13979 => X"88",  -- 136
        13980 => X"88",  -- 136
        13981 => X"8A",  -- 138
        13982 => X"8D",  -- 141
        13983 => X"90",  -- 144
        13984 => X"9D",  -- 157
        13985 => X"A0",  -- 160
        13986 => X"A1",  -- 161
        13987 => X"9E",  -- 158
        13988 => X"99",  -- 153
        13989 => X"95",  -- 149
        13990 => X"96",  -- 150
        13991 => X"98",  -- 152
        13992 => X"90",  -- 144
        13993 => X"8E",  -- 142
        13994 => X"8B",  -- 139
        13995 => X"85",  -- 133
        13996 => X"80",  -- 128
        13997 => X"7D",  -- 125
        13998 => X"7D",  -- 125
        13999 => X"7B",  -- 123
        14000 => X"7F",  -- 127
        14001 => X"90",  -- 144
        14002 => X"95",  -- 149
        14003 => X"83",  -- 131
        14004 => X"75",  -- 117
        14005 => X"7D",  -- 125
        14006 => X"89",  -- 137
        14007 => X"8C",  -- 140
        14008 => X"90",  -- 144
        14009 => X"95",  -- 149
        14010 => X"99",  -- 153
        14011 => X"99",  -- 153
        14012 => X"9B",  -- 155
        14013 => X"9E",  -- 158
        14014 => X"A1",  -- 161
        14015 => X"A1",  -- 161
        14016 => X"A1",  -- 161
        14017 => X"A2",  -- 162
        14018 => X"A6",  -- 166
        14019 => X"AA",  -- 170
        14020 => X"AC",  -- 172
        14021 => X"AB",  -- 171
        14022 => X"A9",  -- 169
        14023 => X"A8",  -- 168
        14024 => X"A4",  -- 164
        14025 => X"9C",  -- 156
        14026 => X"94",  -- 148
        14027 => X"95",  -- 149
        14028 => X"97",  -- 151
        14029 => X"9A",  -- 154
        14030 => X"99",  -- 153
        14031 => X"9B",  -- 155
        14032 => X"98",  -- 152
        14033 => X"93",  -- 147
        14034 => X"8D",  -- 141
        14035 => X"84",  -- 132
        14036 => X"73",  -- 115
        14037 => X"5B",  -- 91
        14038 => X"48",  -- 72
        14039 => X"40",  -- 64
        14040 => X"31",  -- 49
        14041 => X"3F",  -- 63
        14042 => X"58",  -- 88
        14043 => X"75",  -- 117
        14044 => X"88",  -- 136
        14045 => X"8F",  -- 143
        14046 => X"93",  -- 147
        14047 => X"98",  -- 152
        14048 => X"9B",  -- 155
        14049 => X"99",  -- 153
        14050 => X"9A",  -- 154
        14051 => X"98",  -- 152
        14052 => X"97",  -- 151
        14053 => X"9C",  -- 156
        14054 => X"99",  -- 153
        14055 => X"8B",  -- 139
        14056 => X"78",  -- 120
        14057 => X"5C",  -- 92
        14058 => X"55",  -- 85
        14059 => X"6D",  -- 109
        14060 => X"8C",  -- 140
        14061 => X"A2",  -- 162
        14062 => X"AE",  -- 174
        14063 => X"AB",  -- 171
        14064 => X"A8",  -- 168
        14065 => X"A8",  -- 168
        14066 => X"AA",  -- 170
        14067 => X"AC",  -- 172
        14068 => X"B0",  -- 176
        14069 => X"B7",  -- 183
        14070 => X"BF",  -- 191
        14071 => X"C3",  -- 195
        14072 => X"C2",  -- 194
        14073 => X"BC",  -- 188
        14074 => X"C1",  -- 193
        14075 => X"C2",  -- 194
        14076 => X"C1",  -- 193
        14077 => X"B0",  -- 176
        14078 => X"95",  -- 149
        14079 => X"97",  -- 151
        14080 => X"73",  -- 115
        14081 => X"75",  -- 117
        14082 => X"78",  -- 120
        14083 => X"7A",  -- 122
        14084 => X"7A",  -- 122
        14085 => X"75",  -- 117
        14086 => X"70",  -- 112
        14087 => X"6D",  -- 109
        14088 => X"6C",  -- 108
        14089 => X"6A",  -- 106
        14090 => X"69",  -- 105
        14091 => X"6E",  -- 110
        14092 => X"75",  -- 117
        14093 => X"7C",  -- 124
        14094 => X"7C",  -- 124
        14095 => X"7A",  -- 122
        14096 => X"79",  -- 121
        14097 => X"76",  -- 118
        14098 => X"75",  -- 117
        14099 => X"77",  -- 119
        14100 => X"79",  -- 121
        14101 => X"74",  -- 116
        14102 => X"6B",  -- 107
        14103 => X"64",  -- 100
        14104 => X"61",  -- 97
        14105 => X"5F",  -- 95
        14106 => X"59",  -- 89
        14107 => X"4C",  -- 76
        14108 => X"3E",  -- 62
        14109 => X"34",  -- 52
        14110 => X"31",  -- 49
        14111 => X"30",  -- 48
        14112 => X"33",  -- 51
        14113 => X"49",  -- 73
        14114 => X"63",  -- 99
        14115 => X"7B",  -- 123
        14116 => X"90",  -- 144
        14117 => X"99",  -- 153
        14118 => X"8C",  -- 140
        14119 => X"76",  -- 118
        14120 => X"75",  -- 117
        14121 => X"5B",  -- 91
        14122 => X"44",  -- 68
        14123 => X"43",  -- 67
        14124 => X"49",  -- 73
        14125 => X"4A",  -- 74
        14126 => X"48",  -- 72
        14127 => X"49",  -- 73
        14128 => X"4D",  -- 77
        14129 => X"55",  -- 85
        14130 => X"62",  -- 98
        14131 => X"70",  -- 112
        14132 => X"7C",  -- 124
        14133 => X"83",  -- 131
        14134 => X"84",  -- 132
        14135 => X"82",  -- 130
        14136 => X"85",  -- 133
        14137 => X"91",  -- 145
        14138 => X"7B",  -- 123
        14139 => X"61",  -- 97
        14140 => X"4D",  -- 77
        14141 => X"3C",  -- 60
        14142 => X"43",  -- 67
        14143 => X"4D",  -- 77
        14144 => X"56",  -- 86
        14145 => X"51",  -- 81
        14146 => X"6A",  -- 106
        14147 => X"6C",  -- 108
        14148 => X"6A",  -- 106
        14149 => X"6F",  -- 111
        14150 => X"6A",  -- 106
        14151 => X"79",  -- 121
        14152 => X"78",  -- 120
        14153 => X"7D",  -- 125
        14154 => X"74",  -- 116
        14155 => X"63",  -- 99
        14156 => X"45",  -- 69
        14157 => X"40",  -- 64
        14158 => X"33",  -- 51
        14159 => X"30",  -- 48
        14160 => X"1D",  -- 29
        14161 => X"13",  -- 19
        14162 => X"0F",  -- 15
        14163 => X"13",  -- 19
        14164 => X"14",  -- 20
        14165 => X"13",  -- 19
        14166 => X"14",  -- 20
        14167 => X"1C",  -- 28
        14168 => X"12",  -- 18
        14169 => X"12",  -- 18
        14170 => X"13",  -- 19
        14171 => X"0F",  -- 15
        14172 => X"17",  -- 23
        14173 => X"21",  -- 33
        14174 => X"2B",  -- 43
        14175 => X"50",  -- 80
        14176 => X"3B",  -- 59
        14177 => X"40",  -- 64
        14178 => X"32",  -- 50
        14179 => X"20",  -- 32
        14180 => X"1C",  -- 28
        14181 => X"1E",  -- 30
        14182 => X"1B",  -- 27
        14183 => X"1C",  -- 28
        14184 => X"25",  -- 37
        14185 => X"1A",  -- 26
        14186 => X"11",  -- 17
        14187 => X"0D",  -- 13
        14188 => X"0A",  -- 10
        14189 => X"0B",  -- 11
        14190 => X"0C",  -- 12
        14191 => X"12",  -- 18
        14192 => X"19",  -- 25
        14193 => X"15",  -- 21
        14194 => X"17",  -- 23
        14195 => X"19",  -- 25
        14196 => X"19",  -- 25
        14197 => X"24",  -- 36
        14198 => X"35",  -- 53
        14199 => X"3A",  -- 58
        14200 => X"4C",  -- 76
        14201 => X"8B",  -- 139
        14202 => X"8E",  -- 142
        14203 => X"86",  -- 134
        14204 => X"84",  -- 132
        14205 => X"85",  -- 133
        14206 => X"81",  -- 129
        14207 => X"41",  -- 65
        14208 => X"3A",  -- 58
        14209 => X"40",  -- 64
        14210 => X"40",  -- 64
        14211 => X"3A",  -- 58
        14212 => X"3D",  -- 61
        14213 => X"54",  -- 84
        14214 => X"65",  -- 101
        14215 => X"71",  -- 113
        14216 => X"6F",  -- 111
        14217 => X"76",  -- 118
        14218 => X"79",  -- 121
        14219 => X"75",  -- 117
        14220 => X"70",  -- 112
        14221 => X"6A",  -- 106
        14222 => X"5E",  -- 94
        14223 => X"4E",  -- 78
        14224 => X"39",  -- 57
        14225 => X"28",  -- 40
        14226 => X"20",  -- 32
        14227 => X"1D",  -- 29
        14228 => X"16",  -- 22
        14229 => X"21",  -- 33
        14230 => X"2F",  -- 47
        14231 => X"2D",  -- 45
        14232 => X"18",  -- 24
        14233 => X"0D",  -- 13
        14234 => X"05",  -- 5
        14235 => X"17",  -- 23
        14236 => X"4C",  -- 76
        14237 => X"58",  -- 88
        14238 => X"4A",  -- 74
        14239 => X"50",  -- 80
        14240 => X"4E",  -- 78
        14241 => X"47",  -- 71
        14242 => X"45",  -- 69
        14243 => X"4C",  -- 76
        14244 => X"44",  -- 68
        14245 => X"31",  -- 49
        14246 => X"22",  -- 34
        14247 => X"20",  -- 32
        14248 => X"33",  -- 51
        14249 => X"44",  -- 68
        14250 => X"A6",  -- 166
        14251 => X"D1",  -- 209
        14252 => X"A1",  -- 161
        14253 => X"8C",  -- 140
        14254 => X"8A",  -- 138
        14255 => X"7C",  -- 124
        14256 => X"73",  -- 115
        14257 => X"6D",  -- 109
        14258 => X"64",  -- 100
        14259 => X"61",  -- 97
        14260 => X"65",  -- 101
        14261 => X"68",  -- 104
        14262 => X"68",  -- 104
        14263 => X"68",  -- 104
        14264 => X"68",  -- 104
        14265 => X"6B",  -- 107
        14266 => X"6F",  -- 111
        14267 => X"72",  -- 114
        14268 => X"76",  -- 118
        14269 => X"77",  -- 119
        14270 => X"75",  -- 117
        14271 => X"6D",  -- 109
        14272 => X"6D",  -- 109
        14273 => X"6E",  -- 110
        14274 => X"72",  -- 114
        14275 => X"73",  -- 115
        14276 => X"72",  -- 114
        14277 => X"70",  -- 112
        14278 => X"71",  -- 113
        14279 => X"73",  -- 115
        14280 => X"70",  -- 112
        14281 => X"75",  -- 117
        14282 => X"7D",  -- 125
        14283 => X"81",  -- 129
        14284 => X"80",  -- 128
        14285 => X"7D",  -- 125
        14286 => X"7C",  -- 124
        14287 => X"7D",  -- 125
        14288 => X"7F",  -- 127
        14289 => X"7F",  -- 127
        14290 => X"83",  -- 131
        14291 => X"87",  -- 135
        14292 => X"87",  -- 135
        14293 => X"81",  -- 129
        14294 => X"7B",  -- 123
        14295 => X"78",  -- 120
        14296 => X"74",  -- 116
        14297 => X"7D",  -- 125
        14298 => X"86",  -- 134
        14299 => X"8B",  -- 139
        14300 => X"8B",  -- 139
        14301 => X"8B",  -- 139
        14302 => X"91",  -- 145
        14303 => X"98",  -- 152
        14304 => X"9C",  -- 156
        14305 => X"A0",  -- 160
        14306 => X"A1",  -- 161
        14307 => X"9D",  -- 157
        14308 => X"97",  -- 151
        14309 => X"94",  -- 148
        14310 => X"96",  -- 150
        14311 => X"99",  -- 153
        14312 => X"91",  -- 145
        14313 => X"8E",  -- 142
        14314 => X"87",  -- 135
        14315 => X"82",  -- 130
        14316 => X"7F",  -- 127
        14317 => X"7C",  -- 124
        14318 => X"7B",  -- 123
        14319 => X"7B",  -- 123
        14320 => X"7E",  -- 126
        14321 => X"8C",  -- 140
        14322 => X"8F",  -- 143
        14323 => X"7D",  -- 125
        14324 => X"6E",  -- 110
        14325 => X"73",  -- 115
        14326 => X"7C",  -- 124
        14327 => X"7E",  -- 126
        14328 => X"8F",  -- 143
        14329 => X"96",  -- 150
        14330 => X"98",  -- 152
        14331 => X"95",  -- 149
        14332 => X"94",  -- 148
        14333 => X"99",  -- 153
        14334 => X"9D",  -- 157
        14335 => X"9E",  -- 158
        14336 => X"A3",  -- 163
        14337 => X"A6",  -- 166
        14338 => X"A9",  -- 169
        14339 => X"AB",  -- 171
        14340 => X"AD",  -- 173
        14341 => X"AD",  -- 173
        14342 => X"AC",  -- 172
        14343 => X"AB",  -- 171
        14344 => X"AA",  -- 170
        14345 => X"9F",  -- 159
        14346 => X"97",  -- 151
        14347 => X"95",  -- 149
        14348 => X"95",  -- 149
        14349 => X"93",  -- 147
        14350 => X"91",  -- 145
        14351 => X"93",  -- 147
        14352 => X"8D",  -- 141
        14353 => X"89",  -- 137
        14354 => X"87",  -- 135
        14355 => X"80",  -- 128
        14356 => X"71",  -- 113
        14357 => X"54",  -- 84
        14358 => X"39",  -- 57
        14359 => X"2C",  -- 44
        14360 => X"35",  -- 53
        14361 => X"43",  -- 67
        14362 => X"5D",  -- 93
        14363 => X"79",  -- 121
        14364 => X"8C",  -- 140
        14365 => X"93",  -- 147
        14366 => X"95",  -- 149
        14367 => X"97",  -- 151
        14368 => X"98",  -- 152
        14369 => X"95",  -- 149
        14370 => X"97",  -- 151
        14371 => X"94",  -- 148
        14372 => X"92",  -- 146
        14373 => X"98",  -- 152
        14374 => X"95",  -- 149
        14375 => X"86",  -- 134
        14376 => X"6C",  -- 108
        14377 => X"51",  -- 81
        14378 => X"4D",  -- 77
        14379 => X"6A",  -- 106
        14380 => X"8B",  -- 139
        14381 => X"A2",  -- 162
        14382 => X"B0",  -- 176
        14383 => X"B1",  -- 177
        14384 => X"B0",  -- 176
        14385 => X"AD",  -- 173
        14386 => X"AA",  -- 170
        14387 => X"A9",  -- 169
        14388 => X"AE",  -- 174
        14389 => X"B6",  -- 182
        14390 => X"BE",  -- 190
        14391 => X"C2",  -- 194
        14392 => X"C1",  -- 193
        14393 => X"BD",  -- 189
        14394 => X"C3",  -- 195
        14395 => X"BE",  -- 190
        14396 => X"B4",  -- 180
        14397 => X"9D",  -- 157
        14398 => X"8A",  -- 138
        14399 => X"99",  -- 153
        14400 => X"7C",  -- 124
        14401 => X"7C",  -- 124
        14402 => X"7E",  -- 126
        14403 => X"7F",  -- 127
        14404 => X"7E",  -- 126
        14405 => X"79",  -- 121
        14406 => X"73",  -- 115
        14407 => X"6E",  -- 110
        14408 => X"6E",  -- 110
        14409 => X"6B",  -- 107
        14410 => X"67",  -- 103
        14411 => X"69",  -- 105
        14412 => X"6F",  -- 111
        14413 => X"74",  -- 116
        14414 => X"78",  -- 120
        14415 => X"7A",  -- 122
        14416 => X"75",  -- 117
        14417 => X"73",  -- 115
        14418 => X"74",  -- 116
        14419 => X"77",  -- 119
        14420 => X"73",  -- 115
        14421 => X"63",  -- 99
        14422 => X"4C",  -- 76
        14423 => X"3D",  -- 61
        14424 => X"46",  -- 70
        14425 => X"43",  -- 67
        14426 => X"3C",  -- 60
        14427 => X"31",  -- 49
        14428 => X"24",  -- 36
        14429 => X"1B",  -- 27
        14430 => X"19",  -- 25
        14431 => X"1A",  -- 26
        14432 => X"11",  -- 17
        14433 => X"13",  -- 19
        14434 => X"0F",  -- 15
        14435 => X"0F",  -- 15
        14436 => X"20",  -- 32
        14437 => X"4B",  -- 75
        14438 => X"7A",  -- 122
        14439 => X"96",  -- 150
        14440 => X"7B",  -- 123
        14441 => X"5E",  -- 94
        14442 => X"34",  -- 52
        14443 => X"13",  -- 19
        14444 => X"0A",  -- 10
        14445 => X"0E",  -- 14
        14446 => X"0F",  -- 15
        14447 => X"0E",  -- 14
        14448 => X"17",  -- 23
        14449 => X"1D",  -- 29
        14450 => X"24",  -- 36
        14451 => X"32",  -- 50
        14452 => X"46",  -- 70
        14453 => X"5D",  -- 93
        14454 => X"76",  -- 118
        14455 => X"84",  -- 132
        14456 => X"92",  -- 146
        14457 => X"90",  -- 144
        14458 => X"68",  -- 104
        14459 => X"50",  -- 80
        14460 => X"56",  -- 86
        14461 => X"58",  -- 88
        14462 => X"60",  -- 96
        14463 => X"66",  -- 102
        14464 => X"7A",  -- 122
        14465 => X"71",  -- 113
        14466 => X"7A",  -- 122
        14467 => X"79",  -- 121
        14468 => X"72",  -- 114
        14469 => X"7A",  -- 122
        14470 => X"7B",  -- 123
        14471 => X"7E",  -- 126
        14472 => X"79",  -- 121
        14473 => X"62",  -- 98
        14474 => X"3F",  -- 63
        14475 => X"30",  -- 48
        14476 => X"19",  -- 25
        14477 => X"21",  -- 33
        14478 => X"0B",  -- 11
        14479 => X"0D",  -- 13
        14480 => X"0D",  -- 13
        14481 => X"0A",  -- 10
        14482 => X"0C",  -- 12
        14483 => X"12",  -- 18
        14484 => X"14",  -- 20
        14485 => X"12",  -- 18
        14486 => X"12",  -- 18
        14487 => X"13",  -- 19
        14488 => X"17",  -- 23
        14489 => X"11",  -- 17
        14490 => X"12",  -- 18
        14491 => X"10",  -- 16
        14492 => X"15",  -- 21
        14493 => X"1A",  -- 26
        14494 => X"1A",  -- 26
        14495 => X"2C",  -- 44
        14496 => X"3B",  -- 59
        14497 => X"3D",  -- 61
        14498 => X"2D",  -- 45
        14499 => X"1A",  -- 26
        14500 => X"16",  -- 22
        14501 => X"1B",  -- 27
        14502 => X"2B",  -- 43
        14503 => X"3C",  -- 60
        14504 => X"4F",  -- 79
        14505 => X"2B",  -- 43
        14506 => X"25",  -- 37
        14507 => X"2E",  -- 46
        14508 => X"2D",  -- 45
        14509 => X"1C",  -- 28
        14510 => X"10",  -- 16
        14511 => X"22",  -- 34
        14512 => X"20",  -- 32
        14513 => X"1B",  -- 27
        14514 => X"1A",  -- 26
        14515 => X"16",  -- 22
        14516 => X"11",  -- 17
        14517 => X"13",  -- 19
        14518 => X"16",  -- 22
        14519 => X"0E",  -- 14
        14520 => X"2A",  -- 42
        14521 => X"63",  -- 99
        14522 => X"72",  -- 114
        14523 => X"83",  -- 131
        14524 => X"95",  -- 149
        14525 => X"8D",  -- 141
        14526 => X"81",  -- 129
        14527 => X"6A",  -- 106
        14528 => X"77",  -- 119
        14529 => X"6D",  -- 109
        14530 => X"53",  -- 83
        14531 => X"3A",  -- 58
        14532 => X"37",  -- 55
        14533 => X"5E",  -- 94
        14534 => X"6C",  -- 108
        14535 => X"79",  -- 121
        14536 => X"7A",  -- 122
        14537 => X"7E",  -- 126
        14538 => X"7D",  -- 125
        14539 => X"72",  -- 114
        14540 => X"5F",  -- 95
        14541 => X"45",  -- 69
        14542 => X"2A",  -- 42
        14543 => X"18",  -- 24
        14544 => X"0F",  -- 15
        14545 => X"07",  -- 7
        14546 => X"06",  -- 6
        14547 => X"13",  -- 19
        14548 => X"1C",  -- 28
        14549 => X"20",  -- 32
        14550 => X"15",  -- 21
        14551 => X"04",  -- 4
        14552 => X"14",  -- 20
        14553 => X"21",  -- 33
        14554 => X"2C",  -- 44
        14555 => X"3A",  -- 58
        14556 => X"4C",  -- 76
        14557 => X"48",  -- 72
        14558 => X"46",  -- 70
        14559 => X"54",  -- 84
        14560 => X"46",  -- 70
        14561 => X"4F",  -- 79
        14562 => X"57",  -- 87
        14563 => X"50",  -- 80
        14564 => X"45",  -- 69
        14565 => X"3F",  -- 63
        14566 => X"41",  -- 65
        14567 => X"44",  -- 68
        14568 => X"28",  -- 40
        14569 => X"1F",  -- 31
        14570 => X"6C",  -- 108
        14571 => X"AD",  -- 173
        14572 => X"AF",  -- 175
        14573 => X"9A",  -- 154
        14574 => X"78",  -- 120
        14575 => X"6C",  -- 108
        14576 => X"77",  -- 119
        14577 => X"71",  -- 113
        14578 => X"69",  -- 105
        14579 => X"67",  -- 103
        14580 => X"6B",  -- 107
        14581 => X"70",  -- 112
        14582 => X"72",  -- 114
        14583 => X"72",  -- 114
        14584 => X"6C",  -- 108
        14585 => X"6E",  -- 110
        14586 => X"6C",  -- 108
        14587 => X"69",  -- 105
        14588 => X"6A",  -- 106
        14589 => X"6F",  -- 111
        14590 => X"72",  -- 114
        14591 => X"70",  -- 112
        14592 => X"76",  -- 118
        14593 => X"77",  -- 119
        14594 => X"79",  -- 121
        14595 => X"78",  -- 120
        14596 => X"71",  -- 113
        14597 => X"6B",  -- 107
        14598 => X"6C",  -- 108
        14599 => X"71",  -- 113
        14600 => X"72",  -- 114
        14601 => X"75",  -- 117
        14602 => X"7A",  -- 122
        14603 => X"7C",  -- 124
        14604 => X"7A",  -- 122
        14605 => X"77",  -- 119
        14606 => X"7A",  -- 122
        14607 => X"80",  -- 128
        14608 => X"85",  -- 133
        14609 => X"82",  -- 130
        14610 => X"82",  -- 130
        14611 => X"84",  -- 132
        14612 => X"85",  -- 133
        14613 => X"83",  -- 131
        14614 => X"80",  -- 128
        14615 => X"7C",  -- 124
        14616 => X"73",  -- 115
        14617 => X"7B",  -- 123
        14618 => X"85",  -- 133
        14619 => X"8D",  -- 141
        14620 => X"8F",  -- 143
        14621 => X"8F",  -- 143
        14622 => X"95",  -- 149
        14623 => X"9C",  -- 156
        14624 => X"99",  -- 153
        14625 => X"9D",  -- 157
        14626 => X"9D",  -- 157
        14627 => X"9A",  -- 154
        14628 => X"94",  -- 148
        14629 => X"90",  -- 144
        14630 => X"90",  -- 144
        14631 => X"92",  -- 146
        14632 => X"8F",  -- 143
        14633 => X"8A",  -- 138
        14634 => X"83",  -- 131
        14635 => X"80",  -- 128
        14636 => X"81",  -- 129
        14637 => X"82",  -- 130
        14638 => X"82",  -- 130
        14639 => X"81",  -- 129
        14640 => X"87",  -- 135
        14641 => X"83",  -- 131
        14642 => X"83",  -- 131
        14643 => X"80",  -- 128
        14644 => X"70",  -- 112
        14645 => X"60",  -- 96
        14646 => X"66",  -- 102
        14647 => X"78",  -- 120
        14648 => X"8D",  -- 141
        14649 => X"95",  -- 149
        14650 => X"99",  -- 153
        14651 => X"93",  -- 147
        14652 => X"92",  -- 146
        14653 => X"97",  -- 151
        14654 => X"9C",  -- 156
        14655 => X"9C",  -- 156
        14656 => X"A1",  -- 161
        14657 => X"A6",  -- 166
        14658 => X"AB",  -- 171
        14659 => X"AC",  -- 172
        14660 => X"AE",  -- 174
        14661 => X"B1",  -- 177
        14662 => X"B0",  -- 176
        14663 => X"AF",  -- 175
        14664 => X"AC",  -- 172
        14665 => X"A1",  -- 161
        14666 => X"97",  -- 151
        14667 => X"94",  -- 148
        14668 => X"8E",  -- 142
        14669 => X"86",  -- 134
        14670 => X"83",  -- 131
        14671 => X"85",  -- 133
        14672 => X"86",  -- 134
        14673 => X"8A",  -- 138
        14674 => X"8B",  -- 139
        14675 => X"80",  -- 128
        14676 => X"67",  -- 103
        14677 => X"4A",  -- 74
        14678 => X"35",  -- 53
        14679 => X"2E",  -- 46
        14680 => X"39",  -- 57
        14681 => X"44",  -- 68
        14682 => X"57",  -- 87
        14683 => X"71",  -- 113
        14684 => X"84",  -- 132
        14685 => X"8E",  -- 142
        14686 => X"94",  -- 148
        14687 => X"98",  -- 152
        14688 => X"91",  -- 145
        14689 => X"90",  -- 144
        14690 => X"93",  -- 147
        14691 => X"92",  -- 146
        14692 => X"90",  -- 144
        14693 => X"95",  -- 149
        14694 => X"90",  -- 144
        14695 => X"81",  -- 129
        14696 => X"5F",  -- 95
        14697 => X"4B",  -- 75
        14698 => X"4F",  -- 79
        14699 => X"71",  -- 113
        14700 => X"91",  -- 145
        14701 => X"A1",  -- 161
        14702 => X"AA",  -- 170
        14703 => X"AA",  -- 170
        14704 => X"B6",  -- 182
        14705 => X"B2",  -- 178
        14706 => X"AF",  -- 175
        14707 => X"AD",  -- 173
        14708 => X"AE",  -- 174
        14709 => X"B4",  -- 180
        14710 => X"BB",  -- 187
        14711 => X"C0",  -- 192
        14712 => X"BB",  -- 187
        14713 => X"B9",  -- 185
        14714 => X"BE",  -- 190
        14715 => X"B3",  -- 179
        14716 => X"A3",  -- 163
        14717 => X"90",  -- 144
        14718 => X"86",  -- 134
        14719 => X"9E",  -- 158
        14720 => X"88",  -- 136
        14721 => X"87",  -- 135
        14722 => X"86",  -- 134
        14723 => X"86",  -- 134
        14724 => X"85",  -- 133
        14725 => X"81",  -- 129
        14726 => X"7C",  -- 124
        14727 => X"78",  -- 120
        14728 => X"72",  -- 114
        14729 => X"6F",  -- 111
        14730 => X"6C",  -- 108
        14731 => X"6B",  -- 107
        14732 => X"6C",  -- 108
        14733 => X"72",  -- 114
        14734 => X"76",  -- 118
        14735 => X"79",  -- 121
        14736 => X"76",  -- 118
        14737 => X"70",  -- 112
        14738 => X"6D",  -- 109
        14739 => X"69",  -- 105
        14740 => X"5C",  -- 92
        14741 => X"46",  -- 70
        14742 => X"30",  -- 48
        14743 => X"24",  -- 36
        14744 => X"3A",  -- 58
        14745 => X"3B",  -- 59
        14746 => X"3D",  -- 61
        14747 => X"39",  -- 57
        14748 => X"34",  -- 52
        14749 => X"33",  -- 51
        14750 => X"35",  -- 53
        14751 => X"37",  -- 55
        14752 => X"35",  -- 53
        14753 => X"37",  -- 55
        14754 => X"30",  -- 48
        14755 => X"20",  -- 32
        14756 => X"0D",  -- 13
        14757 => X"06",  -- 6
        14758 => X"0B",  -- 11
        14759 => X"13",  -- 19
        14760 => X"56",  -- 86
        14761 => X"59",  -- 89
        14762 => X"40",  -- 64
        14763 => X"16",  -- 22
        14764 => X"05",  -- 5
        14765 => X"0F",  -- 15
        14766 => X"0F",  -- 15
        14767 => X"02",  -- 2
        14768 => X"05",  -- 5
        14769 => X"06",  -- 6
        14770 => X"06",  -- 6
        14771 => X"0C",  -- 12
        14772 => X"1D",  -- 29
        14773 => X"3A",  -- 58
        14774 => X"5D",  -- 93
        14775 => X"76",  -- 118
        14776 => X"86",  -- 134
        14777 => X"84",  -- 132
        14778 => X"5E",  -- 94
        14779 => X"59",  -- 89
        14780 => X"7B",  -- 123
        14781 => X"8B",  -- 139
        14782 => X"8F",  -- 143
        14783 => X"8B",  -- 139
        14784 => X"83",  -- 131
        14785 => X"7D",  -- 125
        14786 => X"79",  -- 121
        14787 => X"7A",  -- 122
        14788 => X"77",  -- 119
        14789 => X"7C",  -- 124
        14790 => X"7E",  -- 126
        14791 => X"66",  -- 102
        14792 => X"52",  -- 82
        14793 => X"32",  -- 50
        14794 => X"1F",  -- 31
        14795 => X"15",  -- 21
        14796 => X"16",  -- 22
        14797 => X"1E",  -- 30
        14798 => X"0E",  -- 14
        14799 => X"12",  -- 18
        14800 => X"1D",  -- 29
        14801 => X"22",  -- 34
        14802 => X"26",  -- 38
        14803 => X"26",  -- 38
        14804 => X"23",  -- 35
        14805 => X"24",  -- 36
        14806 => X"26",  -- 38
        14807 => X"27",  -- 39
        14808 => X"31",  -- 49
        14809 => X"22",  -- 34
        14810 => X"22",  -- 34
        14811 => X"18",  -- 24
        14812 => X"0E",  -- 14
        14813 => X"0E",  -- 14
        14814 => X"08",  -- 8
        14815 => X"08",  -- 8
        14816 => X"1E",  -- 30
        14817 => X"22",  -- 34
        14818 => X"20",  -- 32
        14819 => X"1D",  -- 29
        14820 => X"22",  -- 34
        14821 => X"2B",  -- 43
        14822 => X"42",  -- 66
        14823 => X"60",  -- 96
        14824 => X"74",  -- 116
        14825 => X"56",  -- 86
        14826 => X"5A",  -- 90
        14827 => X"65",  -- 101
        14828 => X"67",  -- 103
        14829 => X"5C",  -- 92
        14830 => X"4A",  -- 74
        14831 => X"57",  -- 87
        14832 => X"51",  -- 81
        14833 => X"45",  -- 69
        14834 => X"38",  -- 56
        14835 => X"2A",  -- 42
        14836 => X"27",  -- 39
        14837 => X"2F",  -- 47
        14838 => X"2A",  -- 42
        14839 => X"16",  -- 22
        14840 => X"17",  -- 23
        14841 => X"28",  -- 40
        14842 => X"3C",  -- 60
        14843 => X"5D",  -- 93
        14844 => X"7A",  -- 122
        14845 => X"7E",  -- 126
        14846 => X"7F",  -- 127
        14847 => X"86",  -- 134
        14848 => X"92",  -- 146
        14849 => X"83",  -- 131
        14850 => X"6B",  -- 107
        14851 => X"50",  -- 80
        14852 => X"43",  -- 67
        14853 => X"62",  -- 98
        14854 => X"63",  -- 99
        14855 => X"73",  -- 115
        14856 => X"79",  -- 121
        14857 => X"76",  -- 118
        14858 => X"6D",  -- 109
        14859 => X"5A",  -- 90
        14860 => X"3F",  -- 63
        14861 => X"20",  -- 32
        14862 => X"0B",  -- 11
        14863 => X"04",  -- 4
        14864 => X"03",  -- 3
        14865 => X"0C",  -- 12
        14866 => X"10",  -- 16
        14867 => X"0B",  -- 11
        14868 => X"07",  -- 7
        14869 => X"07",  -- 7
        14870 => X"12",  -- 18
        14871 => X"26",  -- 38
        14872 => X"24",  -- 36
        14873 => X"2E",  -- 46
        14874 => X"3C",  -- 60
        14875 => X"4A",  -- 74
        14876 => X"53",  -- 83
        14877 => X"59",  -- 89
        14878 => X"5D",  -- 93
        14879 => X"61",  -- 97
        14880 => X"51",  -- 81
        14881 => X"52",  -- 82
        14882 => X"54",  -- 84
        14883 => X"56",  -- 86
        14884 => X"57",  -- 87
        14885 => X"55",  -- 85
        14886 => X"4C",  -- 76
        14887 => X"41",  -- 65
        14888 => X"4D",  -- 77
        14889 => X"34",  -- 52
        14890 => X"1E",  -- 30
        14891 => X"2C",  -- 44
        14892 => X"8A",  -- 138
        14893 => X"B7",  -- 183
        14894 => X"8A",  -- 138
        14895 => X"90",  -- 144
        14896 => X"70",  -- 112
        14897 => X"6B",  -- 107
        14898 => X"65",  -- 101
        14899 => X"65",  -- 101
        14900 => X"6A",  -- 106
        14901 => X"6F",  -- 111
        14902 => X"70",  -- 112
        14903 => X"6F",  -- 111
        14904 => X"6E",  -- 110
        14905 => X"73",  -- 115
        14906 => X"72",  -- 114
        14907 => X"6D",  -- 109
        14908 => X"6B",  -- 107
        14909 => X"6F",  -- 111
        14910 => X"73",  -- 115
        14911 => X"74",  -- 116
        14912 => X"79",  -- 121
        14913 => X"75",  -- 117
        14914 => X"74",  -- 116
        14915 => X"74",  -- 116
        14916 => X"70",  -- 112
        14917 => X"6D",  -- 109
        14918 => X"71",  -- 113
        14919 => X"78",  -- 120
        14920 => X"77",  -- 119
        14921 => X"76",  -- 118
        14922 => X"79",  -- 121
        14923 => X"7C",  -- 124
        14924 => X"7E",  -- 126
        14925 => X"7D",  -- 125
        14926 => X"80",  -- 128
        14927 => X"86",  -- 134
        14928 => X"84",  -- 132
        14929 => X"81",  -- 129
        14930 => X"7F",  -- 127
        14931 => X"80",  -- 128
        14932 => X"84",  -- 132
        14933 => X"86",  -- 134
        14934 => X"83",  -- 131
        14935 => X"7F",  -- 127
        14936 => X"73",  -- 115
        14937 => X"75",  -- 117
        14938 => X"7D",  -- 125
        14939 => X"89",  -- 137
        14940 => X"90",  -- 144
        14941 => X"92",  -- 146
        14942 => X"94",  -- 148
        14943 => X"98",  -- 152
        14944 => X"92",  -- 146
        14945 => X"96",  -- 150
        14946 => X"98",  -- 152
        14947 => X"97",  -- 151
        14948 => X"93",  -- 147
        14949 => X"90",  -- 144
        14950 => X"8E",  -- 142
        14951 => X"8E",  -- 142
        14952 => X"8E",  -- 142
        14953 => X"86",  -- 134
        14954 => X"7D",  -- 125
        14955 => X"7C",  -- 124
        14956 => X"82",  -- 130
        14957 => X"86",  -- 134
        14958 => X"85",  -- 133
        14959 => X"83",  -- 131
        14960 => X"85",  -- 133
        14961 => X"7F",  -- 127
        14962 => X"7F",  -- 127
        14963 => X"81",  -- 129
        14964 => X"6E",  -- 110
        14965 => X"57",  -- 87
        14966 => X"5B",  -- 91
        14967 => X"74",  -- 116
        14968 => X"86",  -- 134
        14969 => X"91",  -- 145
        14970 => X"97",  -- 151
        14971 => X"92",  -- 146
        14972 => X"90",  -- 144
        14973 => X"96",  -- 150
        14974 => X"9A",  -- 154
        14975 => X"9A",  -- 154
        14976 => X"A0",  -- 160
        14977 => X"A7",  -- 167
        14978 => X"AC",  -- 172
        14979 => X"AC",  -- 172
        14980 => X"AE",  -- 174
        14981 => X"B0",  -- 176
        14982 => X"AF",  -- 175
        14983 => X"AC",  -- 172
        14984 => X"A9",  -- 169
        14985 => X"9E",  -- 158
        14986 => X"98",  -- 152
        14987 => X"94",  -- 148
        14988 => X"8C",  -- 140
        14989 => X"81",  -- 129
        14990 => X"7F",  -- 127
        14991 => X"83",  -- 131
        14992 => X"88",  -- 136
        14993 => X"8A",  -- 138
        14994 => X"8B",  -- 139
        14995 => X"80",  -- 128
        14996 => X"68",  -- 104
        14997 => X"4D",  -- 77
        14998 => X"3B",  -- 59
        14999 => X"36",  -- 54
        15000 => X"35",  -- 53
        15001 => X"3C",  -- 60
        15002 => X"4D",  -- 77
        15003 => X"65",  -- 101
        15004 => X"78",  -- 120
        15005 => X"85",  -- 133
        15006 => X"8D",  -- 141
        15007 => X"93",  -- 147
        15008 => X"8C",  -- 140
        15009 => X"8D",  -- 141
        15010 => X"92",  -- 146
        15011 => X"93",  -- 147
        15012 => X"92",  -- 146
        15013 => X"97",  -- 151
        15014 => X"91",  -- 145
        15015 => X"81",  -- 129
        15016 => X"66",  -- 102
        15017 => X"55",  -- 85
        15018 => X"5F",  -- 95
        15019 => X"82",  -- 130
        15020 => X"9E",  -- 158
        15021 => X"A9",  -- 169
        15022 => X"B0",  -- 176
        15023 => X"B1",  -- 177
        15024 => X"B6",  -- 182
        15025 => X"B5",  -- 181
        15026 => X"B5",  -- 181
        15027 => X"B3",  -- 179
        15028 => X"B2",  -- 178
        15029 => X"B4",  -- 180
        15030 => X"BA",  -- 186
        15031 => X"BF",  -- 191
        15032 => X"B9",  -- 185
        15033 => X"B8",  -- 184
        15034 => X"B9",  -- 185
        15035 => X"AA",  -- 170
        15036 => X"9B",  -- 155
        15037 => X"91",  -- 145
        15038 => X"92",  -- 146
        15039 => X"AE",  -- 174
        15040 => X"91",  -- 145
        15041 => X"8F",  -- 143
        15042 => X"8C",  -- 140
        15043 => X"8A",  -- 138
        15044 => X"89",  -- 137
        15045 => X"86",  -- 134
        15046 => X"80",  -- 128
        15047 => X"7B",  -- 123
        15048 => X"79",  -- 121
        15049 => X"77",  -- 119
        15050 => X"74",  -- 116
        15051 => X"72",  -- 114
        15052 => X"71",  -- 113
        15053 => X"74",  -- 116
        15054 => X"79",  -- 121
        15055 => X"7C",  -- 124
        15056 => X"7B",  -- 123
        15057 => X"73",  -- 115
        15058 => X"66",  -- 102
        15059 => X"5B",  -- 91
        15060 => X"4A",  -- 74
        15061 => X"36",  -- 54
        15062 => X"29",  -- 41
        15063 => X"26",  -- 38
        15064 => X"26",  -- 38
        15065 => X"2C",  -- 44
        15066 => X"32",  -- 50
        15067 => X"34",  -- 52
        15068 => X"33",  -- 51
        15069 => X"34",  -- 52
        15070 => X"39",  -- 57
        15071 => X"3D",  -- 61
        15072 => X"44",  -- 68
        15073 => X"39",  -- 57
        15074 => X"33",  -- 51
        15075 => X"40",  -- 64
        15076 => X"4D",  -- 77
        15077 => X"47",  -- 71
        15078 => X"30",  -- 48
        15079 => X"1C",  -- 28
        15080 => X"05",  -- 5
        15081 => X"11",  -- 17
        15082 => X"1C",  -- 28
        15083 => X"1F",  -- 31
        15084 => X"15",  -- 21
        15085 => X"0C",  -- 12
        15086 => X"08",  -- 8
        15087 => X"0A",  -- 10
        15088 => X"08",  -- 8
        15089 => X"0C",  -- 12
        15090 => X"12",  -- 18
        15091 => X"17",  -- 23
        15092 => X"1F",  -- 31
        15093 => X"32",  -- 50
        15094 => X"4A",  -- 74
        15095 => X"5C",  -- 92
        15096 => X"7C",  -- 124
        15097 => X"82",  -- 130
        15098 => X"63",  -- 99
        15099 => X"64",  -- 100
        15100 => X"89",  -- 137
        15101 => X"91",  -- 145
        15102 => X"87",  -- 135
        15103 => X"7D",  -- 125
        15104 => X"79",  -- 121
        15105 => X"79",  -- 121
        15106 => X"6E",  -- 110
        15107 => X"78",  -- 120
        15108 => X"76",  -- 118
        15109 => X"6E",  -- 110
        15110 => X"67",  -- 103
        15111 => X"35",  -- 53
        15112 => X"22",  -- 34
        15113 => X"1A",  -- 26
        15114 => X"34",  -- 52
        15115 => X"2B",  -- 43
        15116 => X"2B",  -- 43
        15117 => X"1E",  -- 30
        15118 => X"24",  -- 36
        15119 => X"3B",  -- 59
        15120 => X"57",  -- 87
        15121 => X"67",  -- 103
        15122 => X"72",  -- 114
        15123 => X"6E",  -- 110
        15124 => X"65",  -- 101
        15125 => X"60",  -- 96
        15126 => X"5D",  -- 93
        15127 => X"59",  -- 89
        15128 => X"64",  -- 100
        15129 => X"51",  -- 81
        15130 => X"50",  -- 80
        15131 => X"39",  -- 57
        15132 => X"1D",  -- 29
        15133 => X"1A",  -- 26
        15134 => X"16",  -- 22
        15135 => X"11",  -- 17
        15136 => X"0A",  -- 10
        15137 => X"13",  -- 19
        15138 => X"1D",  -- 29
        15139 => X"27",  -- 39
        15140 => X"32",  -- 50
        15141 => X"3A",  -- 58
        15142 => X"4E",  -- 78
        15143 => X"6C",  -- 108
        15144 => X"77",  -- 119
        15145 => X"72",  -- 114
        15146 => X"81",  -- 129
        15147 => X"7C",  -- 124
        15148 => X"86",  -- 134
        15149 => X"95",  -- 149
        15150 => X"85",  -- 133
        15151 => X"81",  -- 129
        15152 => X"85",  -- 133
        15153 => X"78",  -- 120
        15154 => X"68",  -- 104
        15155 => X"5A",  -- 90
        15156 => X"5C",  -- 92
        15157 => X"67",  -- 103
        15158 => X"5A",  -- 90
        15159 => X"3A",  -- 58
        15160 => X"18",  -- 24
        15161 => X"09",  -- 9
        15162 => X"16",  -- 22
        15163 => X"2D",  -- 45
        15164 => X"4A",  -- 74
        15165 => X"67",  -- 103
        15166 => X"7A",  -- 122
        15167 => X"8A",  -- 138
        15168 => X"8C",  -- 140
        15169 => X"86",  -- 134
        15170 => X"80",  -- 128
        15171 => X"77",  -- 119
        15172 => X"64",  -- 100
        15173 => X"75",  -- 117
        15174 => X"6B",  -- 107
        15175 => X"7B",  -- 123
        15176 => X"73",  -- 115
        15177 => X"67",  -- 103
        15178 => X"56",  -- 86
        15179 => X"42",  -- 66
        15180 => X"28",  -- 40
        15181 => X"11",  -- 17
        15182 => X"09",  -- 9
        15183 => X"0E",  -- 14
        15184 => X"0E",  -- 14
        15185 => X"0E",  -- 14
        15186 => X"04",  -- 4
        15187 => X"0C",  -- 12
        15188 => X"2B",  -- 43
        15189 => X"39",  -- 57
        15190 => X"35",  -- 53
        15191 => X"39",  -- 57
        15192 => X"3F",  -- 63
        15193 => X"49",  -- 73
        15194 => X"58",  -- 88
        15195 => X"5C",  -- 92
        15196 => X"57",  -- 87
        15197 => X"5A",  -- 90
        15198 => X"5D",  -- 93
        15199 => X"5A",  -- 90
        15200 => X"5B",  -- 91
        15201 => X"55",  -- 85
        15202 => X"50",  -- 80
        15203 => X"4E",  -- 78
        15204 => X"50",  -- 80
        15205 => X"51",  -- 81
        15206 => X"52",  -- 82
        15207 => X"52",  -- 82
        15208 => X"37",  -- 55
        15209 => X"3C",  -- 60
        15210 => X"24",  -- 36
        15211 => X"09",  -- 9
        15212 => X"51",  -- 81
        15213 => X"A4",  -- 164
        15214 => X"88",  -- 136
        15215 => X"77",  -- 119
        15216 => X"77",  -- 119
        15217 => X"71",  -- 113
        15218 => X"6E",  -- 110
        15219 => X"6E",  -- 110
        15220 => X"73",  -- 115
        15221 => X"77",  -- 119
        15222 => X"76",  -- 118
        15223 => X"75",  -- 117
        15224 => X"67",  -- 103
        15225 => X"70",  -- 112
        15226 => X"75",  -- 117
        15227 => X"74",  -- 116
        15228 => X"6F",  -- 111
        15229 => X"6F",  -- 111
        15230 => X"70",  -- 112
        15231 => X"71",  -- 113
        15232 => X"71",  -- 113
        15233 => X"6A",  -- 106
        15234 => X"67",  -- 103
        15235 => X"69",  -- 105
        15236 => X"6C",  -- 108
        15237 => X"6F",  -- 111
        15238 => X"75",  -- 117
        15239 => X"7D",  -- 125
        15240 => X"7E",  -- 126
        15241 => X"7C",  -- 124
        15242 => X"80",  -- 128
        15243 => X"89",  -- 137
        15244 => X"8F",  -- 143
        15245 => X"8E",  -- 142
        15246 => X"8F",  -- 143
        15247 => X"91",  -- 145
        15248 => X"83",  -- 131
        15249 => X"81",  -- 129
        15250 => X"80",  -- 128
        15251 => X"83",  -- 131
        15252 => X"89",  -- 137
        15253 => X"8D",  -- 141
        15254 => X"8A",  -- 138
        15255 => X"86",  -- 134
        15256 => X"74",  -- 116
        15257 => X"71",  -- 113
        15258 => X"77",  -- 119
        15259 => X"86",  -- 134
        15260 => X"93",  -- 147
        15261 => X"96",  -- 150
        15262 => X"95",  -- 149
        15263 => X"94",  -- 148
        15264 => X"8C",  -- 140
        15265 => X"8F",  -- 143
        15266 => X"93",  -- 147
        15267 => X"95",  -- 149
        15268 => X"95",  -- 149
        15269 => X"93",  -- 147
        15270 => X"90",  -- 144
        15271 => X"8F",  -- 143
        15272 => X"8D",  -- 141
        15273 => X"84",  -- 132
        15274 => X"79",  -- 121
        15275 => X"79",  -- 121
        15276 => X"7F",  -- 127
        15277 => X"84",  -- 132
        15278 => X"82",  -- 130
        15279 => X"7E",  -- 126
        15280 => X"7B",  -- 123
        15281 => X"80",  -- 128
        15282 => X"84",  -- 132
        15283 => X"7C",  -- 124
        15284 => X"67",  -- 103
        15285 => X"58",  -- 88
        15286 => X"5F",  -- 95
        15287 => X"70",  -- 112
        15288 => X"7D",  -- 125
        15289 => X"8C",  -- 140
        15290 => X"93",  -- 147
        15291 => X"90",  -- 144
        15292 => X"8F",  -- 143
        15293 => X"95",  -- 149
        15294 => X"98",  -- 152
        15295 => X"96",  -- 150
        15296 => X"A1",  -- 161
        15297 => X"A8",  -- 168
        15298 => X"AD",  -- 173
        15299 => X"AC",  -- 172
        15300 => X"AB",  -- 171
        15301 => X"AC",  -- 172
        15302 => X"AA",  -- 170
        15303 => X"A7",  -- 167
        15304 => X"A5",  -- 165
        15305 => X"9D",  -- 157
        15306 => X"98",  -- 152
        15307 => X"98",  -- 152
        15308 => X"8F",  -- 143
        15309 => X"84",  -- 132
        15310 => X"83",  -- 131
        15311 => X"8A",  -- 138
        15312 => X"8A",  -- 138
        15313 => X"85",  -- 133
        15314 => X"83",  -- 131
        15315 => X"7E",  -- 126
        15316 => X"6F",  -- 111
        15317 => X"58",  -- 88
        15318 => X"40",  -- 64
        15319 => X"33",  -- 51
        15320 => X"35",  -- 53
        15321 => X"3D",  -- 61
        15322 => X"4C",  -- 76
        15323 => X"63",  -- 99
        15324 => X"75",  -- 117
        15325 => X"7F",  -- 127
        15326 => X"84",  -- 132
        15327 => X"88",  -- 136
        15328 => X"8B",  -- 139
        15329 => X"8D",  -- 141
        15330 => X"94",  -- 148
        15331 => X"96",  -- 150
        15332 => X"97",  -- 151
        15333 => X"9B",  -- 155
        15334 => X"95",  -- 149
        15335 => X"84",  -- 132
        15336 => X"67",  -- 103
        15337 => X"54",  -- 84
        15338 => X"5D",  -- 93
        15339 => X"7F",  -- 127
        15340 => X"99",  -- 153
        15341 => X"A4",  -- 164
        15342 => X"AC",  -- 172
        15343 => X"B0",  -- 176
        15344 => X"B4",  -- 180
        15345 => X"B7",  -- 183
        15346 => X"B8",  -- 184
        15347 => X"B7",  -- 183
        15348 => X"B5",  -- 181
        15349 => X"B6",  -- 182
        15350 => X"BA",  -- 186
        15351 => X"BD",  -- 189
        15352 => X"C1",  -- 193
        15353 => X"BF",  -- 191
        15354 => X"BC",  -- 188
        15355 => X"A8",  -- 168
        15356 => X"9B",  -- 155
        15357 => X"96",  -- 150
        15358 => X"9A",  -- 154
        15359 => X"B6",  -- 182
        15360 => X"95",  -- 149
        15361 => X"92",  -- 146
        15362 => X"8E",  -- 142
        15363 => X"89",  -- 137
        15364 => X"84",  -- 132
        15365 => X"82",  -- 130
        15366 => X"81",  -- 129
        15367 => X"80",  -- 128
        15368 => X"7C",  -- 124
        15369 => X"78",  -- 120
        15370 => X"74",  -- 116
        15371 => X"72",  -- 114
        15372 => X"75",  -- 117
        15373 => X"7B",  -- 123
        15374 => X"82",  -- 130
        15375 => X"86",  -- 134
        15376 => X"78",  -- 120
        15377 => X"86",  -- 134
        15378 => X"48",  -- 72
        15379 => X"2C",  -- 44
        15380 => X"2B",  -- 43
        15381 => X"38",  -- 56
        15382 => X"3D",  -- 61
        15383 => X"39",  -- 57
        15384 => X"3E",  -- 62
        15385 => X"4A",  -- 74
        15386 => X"4A",  -- 74
        15387 => X"41",  -- 65
        15388 => X"3F",  -- 63
        15389 => X"47",  -- 71
        15390 => X"4A",  -- 74
        15391 => X"44",  -- 68
        15392 => X"44",  -- 68
        15393 => X"47",  -- 71
        15394 => X"4A",  -- 74
        15395 => X"48",  -- 72
        15396 => X"45",  -- 69
        15397 => X"46",  -- 70
        15398 => X"4B",  -- 75
        15399 => X"4D",  -- 77
        15400 => X"3B",  -- 59
        15401 => X"44",  -- 68
        15402 => X"36",  -- 54
        15403 => X"1F",  -- 31
        15404 => X"12",  -- 18
        15405 => X"0C",  -- 12
        15406 => X"0A",  -- 10
        15407 => X"0C",  -- 12
        15408 => X"0D",  -- 13
        15409 => X"17",  -- 23
        15410 => X"16",  -- 22
        15411 => X"11",  -- 17
        15412 => X"1E",  -- 30
        15413 => X"41",  -- 65
        15414 => X"56",  -- 86
        15415 => X"59",  -- 89
        15416 => X"6D",  -- 109
        15417 => X"71",  -- 113
        15418 => X"64",  -- 100
        15419 => X"6B",  -- 107
        15420 => X"86",  -- 134
        15421 => X"88",  -- 136
        15422 => X"79",  -- 121
        15423 => X"7B",  -- 123
        15424 => X"6A",  -- 106
        15425 => X"7F",  -- 127
        15426 => X"75",  -- 117
        15427 => X"7B",  -- 123
        15428 => X"71",  -- 113
        15429 => X"40",  -- 64
        15430 => X"2D",  -- 45
        15431 => X"2E",  -- 46
        15432 => X"3D",  -- 61
        15433 => X"4B",  -- 75
        15434 => X"53",  -- 83
        15435 => X"6B",  -- 107
        15436 => X"64",  -- 100
        15437 => X"6B",  -- 107
        15438 => X"66",  -- 102
        15439 => X"73",  -- 115
        15440 => X"8B",  -- 139
        15441 => X"85",  -- 133
        15442 => X"77",  -- 119
        15443 => X"80",  -- 128
        15444 => X"7C",  -- 124
        15445 => X"84",  -- 132
        15446 => X"7A",  -- 122
        15447 => X"79",  -- 121
        15448 => X"7B",  -- 123
        15449 => X"70",  -- 112
        15450 => X"6A",  -- 106
        15451 => X"68",  -- 104
        15452 => X"59",  -- 89
        15453 => X"3F",  -- 63
        15454 => X"30",  -- 48
        15455 => X"31",  -- 49
        15456 => X"0B",  -- 11
        15457 => X"1D",  -- 29
        15458 => X"39",  -- 57
        15459 => X"45",  -- 69
        15460 => X"52",  -- 82
        15461 => X"5B",  -- 91
        15462 => X"5E",  -- 94
        15463 => X"6F",  -- 111
        15464 => X"78",  -- 120
        15465 => X"82",  -- 130
        15466 => X"77",  -- 119
        15467 => X"75",  -- 117
        15468 => X"7B",  -- 123
        15469 => X"93",  -- 147
        15470 => X"84",  -- 132
        15471 => X"94",  -- 148
        15472 => X"8B",  -- 139
        15473 => X"89",  -- 137
        15474 => X"90",  -- 144
        15475 => X"8E",  -- 142
        15476 => X"8A",  -- 138
        15477 => X"97",  -- 151
        15478 => X"91",  -- 145
        15479 => X"71",  -- 113
        15480 => X"50",  -- 80
        15481 => X"3C",  -- 60
        15482 => X"26",  -- 38
        15483 => X"23",  -- 35
        15484 => X"31",  -- 49
        15485 => X"45",  -- 69
        15486 => X"60",  -- 96
        15487 => X"81",  -- 129
        15488 => X"8C",  -- 140
        15489 => X"83",  -- 131
        15490 => X"89",  -- 137
        15491 => X"75",  -- 117
        15492 => X"82",  -- 130
        15493 => X"79",  -- 121
        15494 => X"70",  -- 112
        15495 => X"70",  -- 112
        15496 => X"75",  -- 117
        15497 => X"60",  -- 96
        15498 => X"35",  -- 53
        15499 => X"1A",  -- 26
        15500 => X"14",  -- 20
        15501 => X"07",  -- 7
        15502 => X"04",  -- 4
        15503 => X"11",  -- 17
        15504 => X"1B",  -- 27
        15505 => X"18",  -- 24
        15506 => X"1C",  -- 28
        15507 => X"2C",  -- 44
        15508 => X"37",  -- 55
        15509 => X"37",  -- 55
        15510 => X"38",  -- 56
        15511 => X"3E",  -- 62
        15512 => X"47",  -- 71
        15513 => X"59",  -- 89
        15514 => X"53",  -- 83
        15515 => X"5F",  -- 95
        15516 => X"65",  -- 101
        15517 => X"55",  -- 85
        15518 => X"54",  -- 84
        15519 => X"57",  -- 87
        15520 => X"53",  -- 83
        15521 => X"48",  -- 72
        15522 => X"4A",  -- 74
        15523 => X"4D",  -- 77
        15524 => X"46",  -- 70
        15525 => X"50",  -- 80
        15526 => X"55",  -- 85
        15527 => X"4A",  -- 74
        15528 => X"4B",  -- 75
        15529 => X"5B",  -- 91
        15530 => X"3B",  -- 59
        15531 => X"2B",  -- 43
        15532 => X"16",  -- 22
        15533 => X"80",  -- 128
        15534 => X"91",  -- 145
        15535 => X"87",  -- 135
        15536 => X"74",  -- 116
        15537 => X"70",  -- 112
        15538 => X"71",  -- 113
        15539 => X"74",  -- 116
        15540 => X"74",  -- 116
        15541 => X"70",  -- 112
        15542 => X"73",  -- 115
        15543 => X"7B",  -- 123
        15544 => X"7F",  -- 127
        15545 => X"79",  -- 121
        15546 => X"72",  -- 114
        15547 => X"6F",  -- 111
        15548 => X"72",  -- 114
        15549 => X"74",  -- 116
        15550 => X"73",  -- 115
        15551 => X"71",  -- 113
        15552 => X"62",  -- 98
        15553 => X"6D",  -- 109
        15554 => X"78",  -- 120
        15555 => X"79",  -- 121
        15556 => X"71",  -- 113
        15557 => X"6D",  -- 109
        15558 => X"71",  -- 113
        15559 => X"79",  -- 121
        15560 => X"80",  -- 128
        15561 => X"86",  -- 134
        15562 => X"8B",  -- 139
        15563 => X"88",  -- 136
        15564 => X"85",  -- 133
        15565 => X"84",  -- 132
        15566 => X"83",  -- 131
        15567 => X"80",  -- 128
        15568 => X"7C",  -- 124
        15569 => X"7F",  -- 127
        15570 => X"80",  -- 128
        15571 => X"81",  -- 129
        15572 => X"88",  -- 136
        15573 => X"8F",  -- 143
        15574 => X"8E",  -- 142
        15575 => X"88",  -- 136
        15576 => X"79",  -- 121
        15577 => X"71",  -- 113
        15578 => X"72",  -- 114
        15579 => X"81",  -- 129
        15580 => X"8F",  -- 143
        15581 => X"94",  -- 148
        15582 => X"99",  -- 153
        15583 => X"9F",  -- 159
        15584 => X"95",  -- 149
        15585 => X"90",  -- 144
        15586 => X"8D",  -- 141
        15587 => X"90",  -- 144
        15588 => X"91",  -- 145
        15589 => X"8E",  -- 142
        15590 => X"8E",  -- 142
        15591 => X"91",  -- 145
        15592 => X"86",  -- 134
        15593 => X"88",  -- 136
        15594 => X"84",  -- 132
        15595 => X"7C",  -- 124
        15596 => X"7A",  -- 122
        15597 => X"7E",  -- 126
        15598 => X"82",  -- 130
        15599 => X"82",  -- 130
        15600 => X"7A",  -- 122
        15601 => X"80",  -- 128
        15602 => X"81",  -- 129
        15603 => X"7E",  -- 126
        15604 => X"72",  -- 114
        15605 => X"60",  -- 96
        15606 => X"61",  -- 97
        15607 => X"75",  -- 117
        15608 => X"7D",  -- 125
        15609 => X"80",  -- 128
        15610 => X"85",  -- 133
        15611 => X"8B",  -- 139
        15612 => X"8F",  -- 143
        15613 => X"92",  -- 146
        15614 => X"96",  -- 150
        15615 => X"9A",  -- 154
        15616 => X"A0",  -- 160
        15617 => X"A7",  -- 167
        15618 => X"A9",  -- 169
        15619 => X"A5",  -- 165
        15620 => X"A8",  -- 168
        15621 => X"B1",  -- 177
        15622 => X"B5",  -- 181
        15623 => X"B2",  -- 178
        15624 => X"AD",  -- 173
        15625 => X"A2",  -- 162
        15626 => X"96",  -- 150
        15627 => X"90",  -- 144
        15628 => X"91",  -- 145
        15629 => X"90",  -- 144
        15630 => X"89",  -- 137
        15631 => X"83",  -- 131
        15632 => X"86",  -- 134
        15633 => X"7F",  -- 127
        15634 => X"83",  -- 131
        15635 => X"8E",  -- 142
        15636 => X"7D",  -- 125
        15637 => X"55",  -- 85
        15638 => X"38",  -- 56
        15639 => X"35",  -- 53
        15640 => X"3C",  -- 60
        15641 => X"46",  -- 70
        15642 => X"51",  -- 81
        15643 => X"5C",  -- 92
        15644 => X"70",  -- 112
        15645 => X"89",  -- 137
        15646 => X"93",  -- 147
        15647 => X"91",  -- 145
        15648 => X"8F",  -- 143
        15649 => X"93",  -- 147
        15650 => X"93",  -- 147
        15651 => X"93",  -- 147
        15652 => X"97",  -- 151
        15653 => X"9A",  -- 154
        15654 => X"93",  -- 147
        15655 => X"88",  -- 136
        15656 => X"71",  -- 113
        15657 => X"6D",  -- 109
        15658 => X"71",  -- 113
        15659 => X"80",  -- 128
        15660 => X"94",  -- 148
        15661 => X"A5",  -- 165
        15662 => X"AB",  -- 171
        15663 => X"AF",  -- 175
        15664 => X"BA",  -- 186
        15665 => X"BA",  -- 186
        15666 => X"BB",  -- 187
        15667 => X"BA",  -- 186
        15668 => X"B4",  -- 180
        15669 => X"B2",  -- 178
        15670 => X"B8",  -- 184
        15671 => X"BF",  -- 191
        15672 => X"C3",  -- 195
        15673 => X"BA",  -- 186
        15674 => X"B2",  -- 178
        15675 => X"AE",  -- 174
        15676 => X"A5",  -- 165
        15677 => X"9E",  -- 158
        15678 => X"A6",  -- 166
        15679 => X"B7",  -- 183
        15680 => X"8D",  -- 141
        15681 => X"8B",  -- 139
        15682 => X"86",  -- 134
        15683 => X"82",  -- 130
        15684 => X"7F",  -- 127
        15685 => X"7D",  -- 125
        15686 => X"7F",  -- 127
        15687 => X"7F",  -- 127
        15688 => X"83",  -- 131
        15689 => X"81",  -- 129
        15690 => X"7F",  -- 127
        15691 => X"7B",  -- 123
        15692 => X"78",  -- 120
        15693 => X"7A",  -- 122
        15694 => X"7F",  -- 127
        15695 => X"81",  -- 129
        15696 => X"82",  -- 130
        15697 => X"85",  -- 133
        15698 => X"37",  -- 55
        15699 => X"18",  -- 24
        15700 => X"28",  -- 40
        15701 => X"48",  -- 72
        15702 => X"4D",  -- 77
        15703 => X"3F",  -- 63
        15704 => X"44",  -- 68
        15705 => X"4B",  -- 75
        15706 => X"4C",  -- 76
        15707 => X"48",  -- 72
        15708 => X"48",  -- 72
        15709 => X"4E",  -- 78
        15710 => X"4F",  -- 79
        15711 => X"4E",  -- 78
        15712 => X"4F",  -- 79
        15713 => X"56",  -- 86
        15714 => X"54",  -- 84
        15715 => X"4D",  -- 77
        15716 => X"4C",  -- 76
        15717 => X"4D",  -- 77
        15718 => X"43",  -- 67
        15719 => X"32",  -- 50
        15720 => X"4C",  -- 76
        15721 => X"52",  -- 82
        15722 => X"4C",  -- 76
        15723 => X"45",  -- 69
        15724 => X"41",  -- 65
        15725 => X"31",  -- 49
        15726 => X"14",  -- 20
        15727 => X"03",  -- 3
        15728 => X"0E",  -- 14
        15729 => X"10",  -- 16
        15730 => X"0C",  -- 12
        15731 => X"0C",  -- 12
        15732 => X"23",  -- 35
        15733 => X"4A",  -- 74
        15734 => X"63",  -- 99
        15735 => X"6B",  -- 107
        15736 => X"75",  -- 117
        15737 => X"76",  -- 118
        15738 => X"71",  -- 113
        15739 => X"6F",  -- 111
        15740 => X"78",  -- 120
        15741 => X"81",  -- 129
        15742 => X"7D",  -- 125
        15743 => X"73",  -- 115
        15744 => X"79",  -- 121
        15745 => X"7A",  -- 122
        15746 => X"65",  -- 101
        15747 => X"5C",  -- 92
        15748 => X"47",  -- 71
        15749 => X"33",  -- 51
        15750 => X"48",  -- 72
        15751 => X"58",  -- 88
        15752 => X"6E",  -- 110
        15753 => X"86",  -- 134
        15754 => X"8D",  -- 141
        15755 => X"92",  -- 146
        15756 => X"81",  -- 129
        15757 => X"88",  -- 136
        15758 => X"83",  -- 131
        15759 => X"85",  -- 133
        15760 => X"87",  -- 135
        15761 => X"92",  -- 146
        15762 => X"8D",  -- 141
        15763 => X"8A",  -- 138
        15764 => X"7B",  -- 123
        15765 => X"84",  -- 132
        15766 => X"83",  -- 131
        15767 => X"86",  -- 134
        15768 => X"8C",  -- 140
        15769 => X"7C",  -- 124
        15770 => X"73",  -- 115
        15771 => X"73",  -- 115
        15772 => X"69",  -- 105
        15773 => X"52",  -- 82
        15774 => X"4B",  -- 75
        15775 => X"56",  -- 86
        15776 => X"29",  -- 41
        15777 => X"3C",  -- 60
        15778 => X"5B",  -- 91
        15779 => X"5B",  -- 91
        15780 => X"5A",  -- 90
        15781 => X"68",  -- 104
        15782 => X"6F",  -- 111
        15783 => X"77",  -- 119
        15784 => X"75",  -- 117
        15785 => X"6D",  -- 109
        15786 => X"53",  -- 83
        15787 => X"4D",  -- 77
        15788 => X"54",  -- 84
        15789 => X"6B",  -- 107
        15790 => X"5D",  -- 93
        15791 => X"6A",  -- 106
        15792 => X"6D",  -- 109
        15793 => X"6D",  -- 109
        15794 => X"74",  -- 116
        15795 => X"77",  -- 119
        15796 => X"77",  -- 119
        15797 => X"86",  -- 134
        15798 => X"8B",  -- 139
        15799 => X"7A",  -- 122
        15800 => X"97",  -- 151
        15801 => X"82",  -- 130
        15802 => X"6F",  -- 111
        15803 => X"6A",  -- 106
        15804 => X"5A",  -- 90
        15805 => X"39",  -- 57
        15806 => X"33",  -- 51
        15807 => X"4A",  -- 74
        15808 => X"71",  -- 113
        15809 => X"7E",  -- 126
        15810 => X"84",  -- 132
        15811 => X"74",  -- 116
        15812 => X"6C",  -- 108
        15813 => X"76",  -- 118
        15814 => X"70",  -- 112
        15815 => X"78",  -- 120
        15816 => X"71",  -- 113
        15817 => X"51",  -- 81
        15818 => X"28",  -- 40
        15819 => X"12",  -- 18
        15820 => X"0D",  -- 13
        15821 => X"0E",  -- 14
        15822 => X"1E",  -- 30
        15823 => X"38",  -- 56
        15824 => X"2B",  -- 43
        15825 => X"2E",  -- 46
        15826 => X"35",  -- 53
        15827 => X"39",  -- 57
        15828 => X"38",  -- 56
        15829 => X"3B",  -- 59
        15830 => X"4C",  -- 76
        15831 => X"5B",  -- 91
        15832 => X"54",  -- 84
        15833 => X"47",  -- 71
        15834 => X"50",  -- 80
        15835 => X"54",  -- 84
        15836 => X"5E",  -- 94
        15837 => X"6E",  -- 110
        15838 => X"53",  -- 83
        15839 => X"61",  -- 97
        15840 => X"5A",  -- 90
        15841 => X"41",  -- 65
        15842 => X"37",  -- 55
        15843 => X"49",  -- 73
        15844 => X"48",  -- 72
        15845 => X"44",  -- 68
        15846 => X"42",  -- 66
        15847 => X"48",  -- 72
        15848 => X"4D",  -- 77
        15849 => X"54",  -- 84
        15850 => X"4E",  -- 78
        15851 => X"31",  -- 49
        15852 => X"0C",  -- 12
        15853 => X"73",  -- 115
        15854 => X"97",  -- 151
        15855 => X"8C",  -- 140
        15856 => X"84",  -- 132
        15857 => X"76",  -- 118
        15858 => X"6B",  -- 107
        15859 => X"6E",  -- 110
        15860 => X"74",  -- 116
        15861 => X"75",  -- 117
        15862 => X"77",  -- 119
        15863 => X"7B",  -- 123
        15864 => X"77",  -- 119
        15865 => X"72",  -- 114
        15866 => X"6F",  -- 111
        15867 => X"73",  -- 115
        15868 => X"79",  -- 121
        15869 => X"79",  -- 121
        15870 => X"70",  -- 112
        15871 => X"67",  -- 103
        15872 => X"76",  -- 118
        15873 => X"77",  -- 119
        15874 => X"78",  -- 120
        15875 => X"75",  -- 117
        15876 => X"73",  -- 115
        15877 => X"75",  -- 117
        15878 => X"7D",  -- 125
        15879 => X"83",  -- 131
        15880 => X"87",  -- 135
        15881 => X"88",  -- 136
        15882 => X"83",  -- 131
        15883 => X"7D",  -- 125
        15884 => X"7B",  -- 123
        15885 => X"7F",  -- 127
        15886 => X"83",  -- 131
        15887 => X"84",  -- 132
        15888 => X"83",  -- 131
        15889 => X"84",  -- 132
        15890 => X"84",  -- 132
        15891 => X"87",  -- 135
        15892 => X"8D",  -- 141
        15893 => X"94",  -- 148
        15894 => X"95",  -- 149
        15895 => X"91",  -- 145
        15896 => X"79",  -- 121
        15897 => X"73",  -- 115
        15898 => X"76",  -- 118
        15899 => X"86",  -- 134
        15900 => X"94",  -- 148
        15901 => X"97",  -- 151
        15902 => X"98",  -- 152
        15903 => X"9C",  -- 156
        15904 => X"99",  -- 153
        15905 => X"97",  -- 151
        15906 => X"97",  -- 151
        15907 => X"9C",  -- 156
        15908 => X"9C",  -- 156
        15909 => X"97",  -- 151
        15910 => X"93",  -- 147
        15911 => X"93",  -- 147
        15912 => X"90",  -- 144
        15913 => X"8F",  -- 143
        15914 => X"8B",  -- 139
        15915 => X"84",  -- 132
        15916 => X"82",  -- 130
        15917 => X"85",  -- 133
        15918 => X"87",  -- 135
        15919 => X"85",  -- 133
        15920 => X"86",  -- 134
        15921 => X"80",  -- 128
        15922 => X"78",  -- 120
        15923 => X"79",  -- 121
        15924 => X"78",  -- 120
        15925 => X"68",  -- 104
        15926 => X"5F",  -- 95
        15927 => X"68",  -- 104
        15928 => X"6F",  -- 111
        15929 => X"77",  -- 119
        15930 => X"83",  -- 131
        15931 => X"8E",  -- 142
        15932 => X"95",  -- 149
        15933 => X"96",  -- 150
        15934 => X"98",  -- 152
        15935 => X"98",  -- 152
        15936 => X"A1",  -- 161
        15937 => X"A7",  -- 167
        15938 => X"A8",  -- 168
        15939 => X"A6",  -- 166
        15940 => X"AB",  -- 171
        15941 => X"B5",  -- 181
        15942 => X"B7",  -- 183
        15943 => X"B4",  -- 180
        15944 => X"A2",  -- 162
        15945 => X"9C",  -- 156
        15946 => X"98",  -- 152
        15947 => X"98",  -- 152
        15948 => X"98",  -- 152
        15949 => X"94",  -- 148
        15950 => X"89",  -- 137
        15951 => X"80",  -- 128
        15952 => X"82",  -- 130
        15953 => X"7E",  -- 126
        15954 => X"83",  -- 131
        15955 => X"88",  -- 136
        15956 => X"76",  -- 118
        15957 => X"53",  -- 83
        15958 => X"3B",  -- 59
        15959 => X"37",  -- 55
        15960 => X"35",  -- 53
        15961 => X"3D",  -- 61
        15962 => X"4B",  -- 75
        15963 => X"60",  -- 96
        15964 => X"78",  -- 120
        15965 => X"8A",  -- 138
        15966 => X"8E",  -- 142
        15967 => X"8A",  -- 138
        15968 => X"8B",  -- 139
        15969 => X"92",  -- 146
        15970 => X"96",  -- 150
        15971 => X"93",  -- 147
        15972 => X"93",  -- 147
        15973 => X"90",  -- 144
        15974 => X"83",  -- 131
        15975 => X"76",  -- 118
        15976 => X"60",  -- 96
        15977 => X"63",  -- 99
        15978 => X"72",  -- 114
        15979 => X"8C",  -- 140
        15980 => X"A2",  -- 162
        15981 => X"AC",  -- 172
        15982 => X"B1",  -- 177
        15983 => X"B2",  -- 178
        15984 => X"B6",  -- 182
        15985 => X"B7",  -- 183
        15986 => X"B8",  -- 184
        15987 => X"B5",  -- 181
        15988 => X"B1",  -- 177
        15989 => X"B2",  -- 178
        15990 => X"B6",  -- 182
        15991 => X"BE",  -- 190
        15992 => X"BD",  -- 189
        15993 => X"B4",  -- 180
        15994 => X"AF",  -- 175
        15995 => X"B1",  -- 177
        15996 => X"AC",  -- 172
        15997 => X"A6",  -- 166
        15998 => X"AC",  -- 172
        15999 => X"BA",  -- 186
        16000 => X"8D",  -- 141
        16001 => X"89",  -- 137
        16002 => X"85",  -- 133
        16003 => X"81",  -- 129
        16004 => X"7F",  -- 127
        16005 => X"7E",  -- 126
        16006 => X"7F",  -- 127
        16007 => X"80",  -- 128
        16008 => X"84",  -- 132
        16009 => X"85",  -- 133
        16010 => X"83",  -- 131
        16011 => X"7E",  -- 126
        16012 => X"78",  -- 120
        16013 => X"77",  -- 119
        16014 => X"7C",  -- 124
        16015 => X"80",  -- 128
        16016 => X"8F",  -- 143
        16017 => X"6D",  -- 109
        16018 => X"17",  -- 23
        16019 => X"1C",  -- 28
        16020 => X"41",  -- 65
        16021 => X"51",  -- 81
        16022 => X"4D",  -- 77
        16023 => X"4B",  -- 75
        16024 => X"48",  -- 72
        16025 => X"49",  -- 73
        16026 => X"4A",  -- 74
        16027 => X"4B",  -- 75
        16028 => X"4C",  -- 76
        16029 => X"4B",  -- 75
        16030 => X"4C",  -- 76
        16031 => X"4E",  -- 78
        16032 => X"46",  -- 70
        16033 => X"4E",  -- 78
        16034 => X"56",  -- 86
        16035 => X"5A",  -- 90
        16036 => X"5C",  -- 92
        16037 => X"5D",  -- 93
        16038 => X"5B",  -- 91
        16039 => X"56",  -- 86
        16040 => X"45",  -- 69
        16041 => X"49",  -- 73
        16042 => X"46",  -- 70
        16043 => X"49",  -- 73
        16044 => X"55",  -- 85
        16045 => X"51",  -- 81
        16046 => X"41",  -- 65
        16047 => X"38",  -- 56
        16048 => X"19",  -- 25
        16049 => X"17",  -- 23
        16050 => X"14",  -- 20
        16051 => X"13",  -- 19
        16052 => X"20",  -- 32
        16053 => X"3B",  -- 59
        16054 => X"59",  -- 89
        16055 => X"6A",  -- 106
        16056 => X"7A",  -- 122
        16057 => X"70",  -- 112
        16058 => X"6C",  -- 108
        16059 => X"68",  -- 104
        16060 => X"64",  -- 100
        16061 => X"68",  -- 104
        16062 => X"6F",  -- 111
        16063 => X"6E",  -- 110
        16064 => X"5B",  -- 91
        16065 => X"58",  -- 88
        16066 => X"55",  -- 85
        16067 => X"5A",  -- 90
        16068 => X"54",  -- 84
        16069 => X"5C",  -- 92
        16070 => X"7E",  -- 126
        16071 => X"8B",  -- 139
        16072 => X"7F",  -- 127
        16073 => X"92",  -- 146
        16074 => X"90",  -- 144
        16075 => X"86",  -- 134
        16076 => X"7C",  -- 124
        16077 => X"89",  -- 137
        16078 => X"85",  -- 133
        16079 => X"7B",  -- 123
        16080 => X"69",  -- 105
        16081 => X"75",  -- 117
        16082 => X"69",  -- 105
        16083 => X"5C",  -- 92
        16084 => X"49",  -- 73
        16085 => X"5A",  -- 90
        16086 => X"61",  -- 97
        16087 => X"68",  -- 104
        16088 => X"6E",  -- 110
        16089 => X"73",  -- 115
        16090 => X"6F",  -- 111
        16091 => X"6C",  -- 108
        16092 => X"69",  -- 105
        16093 => X"5C",  -- 92
        16094 => X"58",  -- 88
        16095 => X"5F",  -- 95
        16096 => X"47",  -- 71
        16097 => X"45",  -- 69
        16098 => X"6C",  -- 108
        16099 => X"80",  -- 128
        16100 => X"6C",  -- 108
        16101 => X"56",  -- 86
        16102 => X"4F",  -- 79
        16103 => X"5A",  -- 90
        16104 => X"47",  -- 71
        16105 => X"3B",  -- 59
        16106 => X"2C",  -- 44
        16107 => X"28",  -- 40
        16108 => X"2C",  -- 44
        16109 => X"34",  -- 52
        16110 => X"23",  -- 35
        16111 => X"2D",  -- 45
        16112 => X"36",  -- 54
        16113 => X"37",  -- 55
        16114 => X"3F",  -- 63
        16115 => X"44",  -- 68
        16116 => X"45",  -- 69
        16117 => X"51",  -- 81
        16118 => X"5E",  -- 94
        16119 => X"5C",  -- 92
        16120 => X"77",  -- 119
        16121 => X"8B",  -- 139
        16122 => X"93",  -- 147
        16123 => X"8C",  -- 140
        16124 => X"7F",  -- 127
        16125 => X"6B",  -- 107
        16126 => X"55",  -- 85
        16127 => X"4C",  -- 76
        16128 => X"5C",  -- 92
        16129 => X"6F",  -- 111
        16130 => X"75",  -- 117
        16131 => X"72",  -- 114
        16132 => X"63",  -- 99
        16133 => X"7C",  -- 124
        16134 => X"70",  -- 112
        16135 => X"73",  -- 115
        16136 => X"65",  -- 101
        16137 => X"33",  -- 51
        16138 => X"11",  -- 17
        16139 => X"10",  -- 16
        16140 => X"1C",  -- 28
        16141 => X"2D",  -- 45
        16142 => X"3C",  -- 60
        16143 => X"43",  -- 67
        16144 => X"39",  -- 57
        16145 => X"35",  -- 53
        16146 => X"37",  -- 55
        16147 => X"39",  -- 57
        16148 => X"3C",  -- 60
        16149 => X"49",  -- 73
        16150 => X"54",  -- 84
        16151 => X"52",  -- 82
        16152 => X"69",  -- 105
        16153 => X"5D",  -- 93
        16154 => X"5B",  -- 91
        16155 => X"52",  -- 82
        16156 => X"44",  -- 68
        16157 => X"5B",  -- 91
        16158 => X"45",  -- 69
        16159 => X"42",  -- 66
        16160 => X"53",  -- 83
        16161 => X"47",  -- 71
        16162 => X"31",  -- 49
        16163 => X"3F",  -- 63
        16164 => X"40",  -- 64
        16165 => X"49",  -- 73
        16166 => X"42",  -- 66
        16167 => X"52",  -- 82
        16168 => X"4F",  -- 79
        16169 => X"45",  -- 69
        16170 => X"59",  -- 89
        16171 => X"37",  -- 55
        16172 => X"0B",  -- 11
        16173 => X"6C",  -- 108
        16174 => X"B1",  -- 177
        16175 => X"9A",  -- 154
        16176 => X"7F",  -- 127
        16177 => X"76",  -- 118
        16178 => X"72",  -- 114
        16179 => X"79",  -- 121
        16180 => X"7D",  -- 125
        16181 => X"79",  -- 121
        16182 => X"75",  -- 117
        16183 => X"76",  -- 118
        16184 => X"71",  -- 113
        16185 => X"72",  -- 114
        16186 => X"74",  -- 116
        16187 => X"77",  -- 119
        16188 => X"7A",  -- 122
        16189 => X"79",  -- 121
        16190 => X"74",  -- 116
        16191 => X"6F",  -- 111
        16192 => X"82",  -- 130
        16193 => X"7B",  -- 123
        16194 => X"75",  -- 117
        16195 => X"72",  -- 114
        16196 => X"75",  -- 117
        16197 => X"7B",  -- 123
        16198 => X"81",  -- 129
        16199 => X"84",  -- 132
        16200 => X"7C",  -- 124
        16201 => X"7F",  -- 127
        16202 => X"80",  -- 128
        16203 => X"80",  -- 128
        16204 => X"85",  -- 133
        16205 => X"8A",  -- 138
        16206 => X"8C",  -- 140
        16207 => X"89",  -- 137
        16208 => X"86",  -- 134
        16209 => X"86",  -- 134
        16210 => X"86",  -- 134
        16211 => X"86",  -- 134
        16212 => X"8B",  -- 139
        16213 => X"91",  -- 145
        16214 => X"93",  -- 147
        16215 => X"90",  -- 144
        16216 => X"84",  -- 132
        16217 => X"7B",  -- 123
        16218 => X"79",  -- 121
        16219 => X"86",  -- 134
        16220 => X"94",  -- 148
        16221 => X"9A",  -- 154
        16222 => X"9B",  -- 155
        16223 => X"9D",  -- 157
        16224 => X"9F",  -- 159
        16225 => X"9E",  -- 158
        16226 => X"9F",  -- 159
        16227 => X"A2",  -- 162
        16228 => X"A2",  -- 162
        16229 => X"9E",  -- 158
        16230 => X"99",  -- 153
        16231 => X"98",  -- 152
        16232 => X"98",  -- 152
        16233 => X"94",  -- 148
        16234 => X"8C",  -- 140
        16235 => X"86",  -- 134
        16236 => X"85",  -- 133
        16237 => X"87",  -- 135
        16238 => X"85",  -- 133
        16239 => X"82",  -- 130
        16240 => X"86",  -- 134
        16241 => X"7E",  -- 126
        16242 => X"74",  -- 116
        16243 => X"75",  -- 117
        16244 => X"79",  -- 121
        16245 => X"6B",  -- 107
        16246 => X"5F",  -- 95
        16247 => X"63",  -- 99
        16248 => X"73",  -- 115
        16249 => X"7E",  -- 126
        16250 => X"8D",  -- 141
        16251 => X"98",  -- 152
        16252 => X"9E",  -- 158
        16253 => X"A0",  -- 160
        16254 => X"A2",  -- 162
        16255 => X"A2",  -- 162
        16256 => X"A0",  -- 160
        16257 => X"A4",  -- 164
        16258 => X"A5",  -- 165
        16259 => X"A6",  -- 166
        16260 => X"AD",  -- 173
        16261 => X"B6",  -- 182
        16262 => X"B6",  -- 182
        16263 => X"B1",  -- 177
        16264 => X"A4",  -- 164
        16265 => X"A0",  -- 160
        16266 => X"9C",  -- 156
        16267 => X"9D",  -- 157
        16268 => X"9B",  -- 155
        16269 => X"96",  -- 150
        16270 => X"8C",  -- 140
        16271 => X"82",  -- 130
        16272 => X"76",  -- 118
        16273 => X"78",  -- 120
        16274 => X"7F",  -- 127
        16275 => X"7E",  -- 126
        16276 => X"6C",  -- 108
        16277 => X"50",  -- 80
        16278 => X"3E",  -- 62
        16279 => X"38",  -- 56
        16280 => X"2D",  -- 45
        16281 => X"2F",  -- 47
        16282 => X"3E",  -- 62
        16283 => X"5A",  -- 90
        16284 => X"74",  -- 116
        16285 => X"81",  -- 129
        16286 => X"83",  -- 131
        16287 => X"83",  -- 131
        16288 => X"8A",  -- 138
        16289 => X"91",  -- 145
        16290 => X"95",  -- 149
        16291 => X"92",  -- 146
        16292 => X"90",  -- 144
        16293 => X"8A",  -- 138
        16294 => X"7D",  -- 125
        16295 => X"6D",  -- 109
        16296 => X"57",  -- 87
        16297 => X"5F",  -- 95
        16298 => X"75",  -- 117
        16299 => X"94",  -- 148
        16300 => X"A7",  -- 167
        16301 => X"AB",  -- 171
        16302 => X"AF",  -- 175
        16303 => X"B4",  -- 180
        16304 => X"B5",  -- 181
        16305 => X"B6",  -- 182
        16306 => X"B6",  -- 182
        16307 => X"B2",  -- 178
        16308 => X"AF",  -- 175
        16309 => X"B2",  -- 178
        16310 => X"B9",  -- 185
        16311 => X"BE",  -- 190
        16312 => X"BD",  -- 189
        16313 => X"B6",  -- 182
        16314 => X"B5",  -- 181
        16315 => X"B9",  -- 185
        16316 => X"B8",  -- 184
        16317 => X"B3",  -- 179
        16318 => X"B6",  -- 182
        16319 => X"C0",  -- 192
        16320 => X"8D",  -- 141
        16321 => X"8B",  -- 139
        16322 => X"86",  -- 134
        16323 => X"83",  -- 131
        16324 => X"7F",  -- 127
        16325 => X"7D",  -- 125
        16326 => X"7C",  -- 124
        16327 => X"7C",  -- 124
        16328 => X"7B",  -- 123
        16329 => X"7E",  -- 126
        16330 => X"7D",  -- 125
        16331 => X"79",  -- 121
        16332 => X"74",  -- 116
        16333 => X"74",  -- 116
        16334 => X"7B",  -- 123
        16335 => X"83",  -- 131
        16336 => X"8E",  -- 142
        16337 => X"72",  -- 114
        16338 => X"2A",  -- 42
        16339 => X"3B",  -- 59
        16340 => X"54",  -- 84
        16341 => X"4F",  -- 79
        16342 => X"49",  -- 73
        16343 => X"53",  -- 83
        16344 => X"49",  -- 73
        16345 => X"45",  -- 69
        16346 => X"45",  -- 69
        16347 => X"49",  -- 73
        16348 => X"48",  -- 72
        16349 => X"3F",  -- 63
        16350 => X"3C",  -- 60
        16351 => X"40",  -- 64
        16352 => X"30",  -- 48
        16353 => X"3C",  -- 60
        16354 => X"53",  -- 83
        16355 => X"61",  -- 97
        16356 => X"59",  -- 89
        16357 => X"4B",  -- 75
        16358 => X"50",  -- 80
        16359 => X"62",  -- 98
        16360 => X"51",  -- 81
        16361 => X"53",  -- 83
        16362 => X"49",  -- 73
        16363 => X"40",  -- 64
        16364 => X"42",  -- 66
        16365 => X"46",  -- 70
        16366 => X"4F",  -- 79
        16367 => X"5C",  -- 92
        16368 => X"55",  -- 85
        16369 => X"4E",  -- 78
        16370 => X"3F",  -- 63
        16371 => X"29",  -- 41
        16372 => X"1C",  -- 28
        16373 => X"2A",  -- 42
        16374 => X"55",  -- 85
        16375 => X"7A",  -- 122
        16376 => X"87",  -- 135
        16377 => X"78",  -- 120
        16378 => X"6A",  -- 106
        16379 => X"69",  -- 105
        16380 => X"67",  -- 103
        16381 => X"59",  -- 89
        16382 => X"57",  -- 87
        16383 => X"63",  -- 99
        16384 => X"4F",  -- 79
        16385 => X"5A",  -- 90
        16386 => X"65",  -- 101
        16387 => X"7A",  -- 122
        16388 => X"8D",  -- 141
        16389 => X"8E",  -- 142
        16390 => X"8B",  -- 139
        16391 => X"88",  -- 136
        16392 => X"70",  -- 112
        16393 => X"6B",  -- 107
        16394 => X"58",  -- 88
        16395 => X"47",  -- 71
        16396 => X"44",  -- 68
        16397 => X"50",  -- 80
        16398 => X"46",  -- 70
        16399 => X"34",  -- 52
        16400 => X"38",  -- 56
        16401 => X"38",  -- 56
        16402 => X"2A",  -- 42
        16403 => X"29",  -- 41
        16404 => X"21",  -- 33
        16405 => X"2D",  -- 45
        16406 => X"2B",  -- 43
        16407 => X"2D",  -- 45
        16408 => X"39",  -- 57
        16409 => X"4D",  -- 77
        16410 => X"4B",  -- 75
        16411 => X"42",  -- 66
        16412 => X"4C",  -- 76
        16413 => X"57",  -- 87
        16414 => X"5C",  -- 92
        16415 => X"5F",  -- 95
        16416 => X"51",  -- 81
        16417 => X"45",  -- 69
        16418 => X"69",  -- 105
        16419 => X"7A",  -- 122
        16420 => X"5E",  -- 94
        16421 => X"43",  -- 67
        16422 => X"30",  -- 48
        16423 => X"28",  -- 40
        16424 => X"24",  -- 36
        16425 => X"1E",  -- 30
        16426 => X"1F",  -- 31
        16427 => X"1F",  -- 31
        16428 => X"1B",  -- 27
        16429 => X"18",  -- 24
        16430 => X"0F",  -- 15
        16431 => X"1A",  -- 26
        16432 => X"14",  -- 20
        16433 => X"15",  -- 21
        16434 => X"1C",  -- 28
        16435 => X"20",  -- 32
        16436 => X"1C",  -- 28
        16437 => X"1E",  -- 30
        16438 => X"29",  -- 41
        16439 => X"32",  -- 50
        16440 => X"3B",  -- 59
        16441 => X"61",  -- 97
        16442 => X"75",  -- 117
        16443 => X"79",  -- 121
        16444 => X"88",  -- 136
        16445 => X"94",  -- 148
        16446 => X"7F",  -- 127
        16447 => X"62",  -- 98
        16448 => X"5A",  -- 90
        16449 => X"58",  -- 88
        16450 => X"61",  -- 97
        16451 => X"6E",  -- 110
        16452 => X"74",  -- 116
        16453 => X"85",  -- 133
        16454 => X"6C",  -- 108
        16455 => X"5B",  -- 91
        16456 => X"49",  -- 73
        16457 => X"28",  -- 40
        16458 => X"1D",  -- 29
        16459 => X"2A",  -- 42
        16460 => X"38",  -- 56
        16461 => X"45",  -- 69
        16462 => X"44",  -- 68
        16463 => X"30",  -- 48
        16464 => X"28",  -- 40
        16465 => X"2D",  -- 45
        16466 => X"3F",  -- 63
        16467 => X"4D",  -- 77
        16468 => X"52",  -- 82
        16469 => X"5B",  -- 91
        16470 => X"52",  -- 82
        16471 => X"37",  -- 55
        16472 => X"4B",  -- 75
        16473 => X"6B",  -- 107
        16474 => X"61",  -- 97
        16475 => X"6C",  -- 108
        16476 => X"4C",  -- 76
        16477 => X"51",  -- 81
        16478 => X"5F",  -- 95
        16479 => X"46",  -- 70
        16480 => X"55",  -- 85
        16481 => X"68",  -- 104
        16482 => X"4E",  -- 78
        16483 => X"3A",  -- 58
        16484 => X"2F",  -- 47
        16485 => X"47",  -- 71
        16486 => X"40",  -- 64
        16487 => X"44",  -- 68
        16488 => X"5A",  -- 90
        16489 => X"48",  -- 72
        16490 => X"59",  -- 89
        16491 => X"40",  -- 64
        16492 => X"17",  -- 23
        16493 => X"5D",  -- 93
        16494 => X"C6",  -- 198
        16495 => X"A4",  -- 164
        16496 => X"7D",  -- 125
        16497 => X"7D",  -- 125
        16498 => X"7F",  -- 127
        16499 => X"7F",  -- 127
        16500 => X"76",  -- 118
        16501 => X"6A",  -- 106
        16502 => X"6A",  -- 106
        16503 => X"71",  -- 113
        16504 => X"71",  -- 113
        16505 => X"75",  -- 117
        16506 => X"77",  -- 119
        16507 => X"74",  -- 116
        16508 => X"70",  -- 112
        16509 => X"72",  -- 114
        16510 => X"7C",  -- 124
        16511 => X"86",  -- 134
        16512 => X"81",  -- 129
        16513 => X"7C",  -- 124
        16514 => X"77",  -- 119
        16515 => X"77",  -- 119
        16516 => X"7B",  -- 123
        16517 => X"7E",  -- 126
        16518 => X"7E",  -- 126
        16519 => X"7D",  -- 125
        16520 => X"7A",  -- 122
        16521 => X"7E",  -- 126
        16522 => X"81",  -- 129
        16523 => X"86",  -- 134
        16524 => X"8D",  -- 141
        16525 => X"95",  -- 149
        16526 => X"94",  -- 148
        16527 => X"8F",  -- 143
        16528 => X"91",  -- 145
        16529 => X"91",  -- 145
        16530 => X"8D",  -- 141
        16531 => X"8C",  -- 140
        16532 => X"8D",  -- 141
        16533 => X"8F",  -- 143
        16534 => X"8F",  -- 143
        16535 => X"8F",  -- 143
        16536 => X"91",  -- 145
        16537 => X"80",  -- 128
        16538 => X"74",  -- 116
        16539 => X"7A",  -- 122
        16540 => X"8C",  -- 140
        16541 => X"97",  -- 151
        16542 => X"9D",  -- 157
        16543 => X"9F",  -- 159
        16544 => X"A1",  -- 161
        16545 => X"A0",  -- 160
        16546 => X"9E",  -- 158
        16547 => X"9E",  -- 158
        16548 => X"9F",  -- 159
        16549 => X"9D",  -- 157
        16550 => X"9C",  -- 156
        16551 => X"9B",  -- 155
        16552 => X"96",  -- 150
        16553 => X"90",  -- 144
        16554 => X"88",  -- 136
        16555 => X"83",  -- 131
        16556 => X"83",  -- 131
        16557 => X"83",  -- 131
        16558 => X"80",  -- 128
        16559 => X"7B",  -- 123
        16560 => X"79",  -- 121
        16561 => X"7B",  -- 123
        16562 => X"79",  -- 121
        16563 => X"78",  -- 120
        16564 => X"72",  -- 114
        16565 => X"61",  -- 97
        16566 => X"5C",  -- 92
        16567 => X"67",  -- 103
        16568 => X"6E",  -- 110
        16569 => X"79",  -- 121
        16570 => X"85",  -- 133
        16571 => X"8D",  -- 141
        16572 => X"93",  -- 147
        16573 => X"98",  -- 152
        16574 => X"9C",  -- 156
        16575 => X"9F",  -- 159
        16576 => X"9E",  -- 158
        16577 => X"A0",  -- 160
        16578 => X"A1",  -- 161
        16579 => X"A4",  -- 164
        16580 => X"AC",  -- 172
        16581 => X"B2",  -- 178
        16582 => X"B0",  -- 176
        16583 => X"AA",  -- 170
        16584 => X"AC",  -- 172
        16585 => X"A5",  -- 165
        16586 => X"9B",  -- 155
        16587 => X"95",  -- 149
        16588 => X"91",  -- 145
        16589 => X"8C",  -- 140
        16590 => X"87",  -- 135
        16591 => X"81",  -- 129
        16592 => X"71",  -- 113
        16593 => X"76",  -- 118
        16594 => X"7C",  -- 124
        16595 => X"7A",  -- 122
        16596 => X"6C",  -- 108
        16597 => X"57",  -- 87
        16598 => X"44",  -- 68
        16599 => X"38",  -- 56
        16600 => X"2A",  -- 42
        16601 => X"2A",  -- 42
        16602 => X"39",  -- 57
        16603 => X"55",  -- 85
        16604 => X"6E",  -- 110
        16605 => X"78",  -- 120
        16606 => X"7F",  -- 127
        16607 => X"88",  -- 136
        16608 => X"91",  -- 145
        16609 => X"95",  -- 149
        16610 => X"95",  -- 149
        16611 => X"95",  -- 149
        16612 => X"97",  -- 151
        16613 => X"95",  -- 149
        16614 => X"85",  -- 133
        16615 => X"74",  -- 116
        16616 => X"60",  -- 96
        16617 => X"69",  -- 105
        16618 => X"7F",  -- 127
        16619 => X"98",  -- 152
        16620 => X"A4",  -- 164
        16621 => X"A5",  -- 165
        16622 => X"AB",  -- 171
        16623 => X"B5",  -- 181
        16624 => X"B7",  -- 183
        16625 => X"B7",  -- 183
        16626 => X"B6",  -- 182
        16627 => X"B1",  -- 177
        16628 => X"B1",  -- 177
        16629 => X"B6",  -- 182
        16630 => X"BD",  -- 189
        16631 => X"C2",  -- 194
        16632 => X"C1",  -- 193
        16633 => X"B8",  -- 184
        16634 => X"B7",  -- 183
        16635 => X"BF",  -- 191
        16636 => X"C0",  -- 192
        16637 => X"B9",  -- 185
        16638 => X"BA",  -- 186
        16639 => X"C2",  -- 194
        16640 => X"83",  -- 131
        16641 => X"83",  -- 131
        16642 => X"82",  -- 130
        16643 => X"80",  -- 128
        16644 => X"7D",  -- 125
        16645 => X"79",  -- 121
        16646 => X"76",  -- 118
        16647 => X"74",  -- 116
        16648 => X"73",  -- 115
        16649 => X"75",  -- 117
        16650 => X"76",  -- 118
        16651 => X"73",  -- 115
        16652 => X"70",  -- 112
        16653 => X"73",  -- 115
        16654 => X"7D",  -- 125
        16655 => X"84",  -- 132
        16656 => X"85",  -- 133
        16657 => X"8D",  -- 141
        16658 => X"50",  -- 80
        16659 => X"40",  -- 64
        16660 => X"47",  -- 71
        16661 => X"51",  -- 81
        16662 => X"52",  -- 82
        16663 => X"4E",  -- 78
        16664 => X"47",  -- 71
        16665 => X"42",  -- 66
        16666 => X"42",  -- 66
        16667 => X"47",  -- 71
        16668 => X"44",  -- 68
        16669 => X"3B",  -- 59
        16670 => X"37",  -- 55
        16671 => X"3A",  -- 58
        16672 => X"46",  -- 70
        16673 => X"58",  -- 88
        16674 => X"68",  -- 104
        16675 => X"65",  -- 101
        16676 => X"52",  -- 82
        16677 => X"44",  -- 68
        16678 => X"43",  -- 67
        16679 => X"4B",  -- 75
        16680 => X"58",  -- 88
        16681 => X"60",  -- 96
        16682 => X"5A",  -- 90
        16683 => X"49",  -- 73
        16684 => X"41",  -- 65
        16685 => X"42",  -- 66
        16686 => X"48",  -- 72
        16687 => X"53",  -- 83
        16688 => X"60",  -- 96
        16689 => X"66",  -- 102
        16690 => X"67",  -- 103
        16691 => X"5C",  -- 92
        16692 => X"49",  -- 73
        16693 => X"41",  -- 65
        16694 => X"51",  -- 81
        16695 => X"66",  -- 102
        16696 => X"85",  -- 133
        16697 => X"8E",  -- 142
        16698 => X"80",  -- 128
        16699 => X"7A",  -- 122
        16700 => X"83",  -- 131
        16701 => X"6B",  -- 107
        16702 => X"4C",  -- 76
        16703 => X"4C",  -- 76
        16704 => X"69",  -- 105
        16705 => X"7C",  -- 124
        16706 => X"84",  -- 132
        16707 => X"8C",  -- 140
        16708 => X"98",  -- 152
        16709 => X"7D",  -- 125
        16710 => X"53",  -- 83
        16711 => X"4F",  -- 79
        16712 => X"3A",  -- 58
        16713 => X"29",  -- 41
        16714 => X"1A",  -- 26
        16715 => X"13",  -- 19
        16716 => X"19",  -- 25
        16717 => X"1A",  -- 26
        16718 => X"17",  -- 23
        16719 => X"10",  -- 16
        16720 => X"15",  -- 21
        16721 => X"12",  -- 18
        16722 => X"10",  -- 16
        16723 => X"23",  -- 35
        16724 => X"1E",  -- 30
        16725 => X"1D",  -- 29
        16726 => X"11",  -- 17
        16727 => X"18",  -- 24
        16728 => X"1D",  -- 29
        16729 => X"21",  -- 33
        16730 => X"15",  -- 21
        16731 => X"13",  -- 19
        16732 => X"28",  -- 40
        16733 => X"38",  -- 56
        16734 => X"47",  -- 71
        16735 => X"61",  -- 97
        16736 => X"4C",  -- 76
        16737 => X"56",  -- 86
        16738 => X"6B",  -- 107
        16739 => X"58",  -- 88
        16740 => X"49",  -- 73
        16741 => X"5E",  -- 94
        16742 => X"53",  -- 83
        16743 => X"2B",  -- 43
        16744 => X"22",  -- 34
        16745 => X"16",  -- 22
        16746 => X"1C",  -- 28
        16747 => X"18",  -- 24
        16748 => X"16",  -- 22
        16749 => X"13",  -- 19
        16750 => X"10",  -- 16
        16751 => X"1A",  -- 26
        16752 => X"11",  -- 17
        16753 => X"15",  -- 21
        16754 => X"1A",  -- 26
        16755 => X"1D",  -- 29
        16756 => X"1B",  -- 27
        16757 => X"16",  -- 22
        16758 => X"19",  -- 25
        16759 => X"23",  -- 35
        16760 => X"2E",  -- 46
        16761 => X"34",  -- 52
        16762 => X"3C",  -- 60
        16763 => X"54",  -- 84
        16764 => X"77",  -- 119
        16765 => X"87",  -- 135
        16766 => X"7C",  -- 124
        16767 => X"73",  -- 115
        16768 => X"55",  -- 85
        16769 => X"3F",  -- 63
        16770 => X"55",  -- 85
        16771 => X"69",  -- 105
        16772 => X"81",  -- 129
        16773 => X"7D",  -- 125
        16774 => X"63",  -- 99
        16775 => X"46",  -- 70
        16776 => X"3B",  -- 59
        16777 => X"3C",  -- 60
        16778 => X"4A",  -- 74
        16779 => X"4C",  -- 76
        16780 => X"40",  -- 64
        16781 => X"3F",  -- 63
        16782 => X"3C",  -- 60
        16783 => X"2A",  -- 42
        16784 => X"30",  -- 48
        16785 => X"38",  -- 56
        16786 => X"4D",  -- 77
        16787 => X"53",  -- 83
        16788 => X"4C",  -- 76
        16789 => X"5B",  -- 91
        16790 => X"68",  -- 104
        16791 => X"58",  -- 88
        16792 => X"60",  -- 96
        16793 => X"78",  -- 120
        16794 => X"73",  -- 115
        16795 => X"8E",  -- 142
        16796 => X"68",  -- 104
        16797 => X"4D",  -- 77
        16798 => X"61",  -- 97
        16799 => X"55",  -- 85
        16800 => X"47",  -- 71
        16801 => X"70",  -- 112
        16802 => X"66",  -- 102
        16803 => X"45",  -- 69
        16804 => X"34",  -- 52
        16805 => X"4A",  -- 74
        16806 => X"49",  -- 73
        16807 => X"49",  -- 73
        16808 => X"60",  -- 96
        16809 => X"5B",  -- 91
        16810 => X"5E",  -- 94
        16811 => X"50",  -- 80
        16812 => X"28",  -- 40
        16813 => X"3D",  -- 61
        16814 => X"BF",  -- 191
        16815 => X"A7",  -- 167
        16816 => X"94",  -- 148
        16817 => X"88",  -- 136
        16818 => X"7C",  -- 124
        16819 => X"72",  -- 114
        16820 => X"67",  -- 103
        16821 => X"60",  -- 96
        16822 => X"67",  -- 103
        16823 => X"74",  -- 116
        16824 => X"72",  -- 114
        16825 => X"70",  -- 112
        16826 => X"6D",  -- 109
        16827 => X"69",  -- 105
        16828 => X"6A",  -- 106
        16829 => X"72",  -- 114
        16830 => X"7E",  -- 126
        16831 => X"88",  -- 136
        16832 => X"81",  -- 129
        16833 => X"7F",  -- 127
        16834 => X"7E",  -- 126
        16835 => X"7F",  -- 127
        16836 => X"81",  -- 129
        16837 => X"81",  -- 129
        16838 => X"80",  -- 128
        16839 => X"7F",  -- 127
        16840 => X"84",  -- 132
        16841 => X"82",  -- 130
        16842 => X"7E",  -- 126
        16843 => X"7B",  -- 123
        16844 => X"81",  -- 129
        16845 => X"8A",  -- 138
        16846 => X"90",  -- 144
        16847 => X"90",  -- 144
        16848 => X"9D",  -- 157
        16849 => X"9C",  -- 156
        16850 => X"99",  -- 153
        16851 => X"98",  -- 152
        16852 => X"98",  -- 152
        16853 => X"96",  -- 150
        16854 => X"96",  -- 150
        16855 => X"95",  -- 149
        16856 => X"8F",  -- 143
        16857 => X"7D",  -- 125
        16858 => X"6E",  -- 110
        16859 => X"73",  -- 115
        16860 => X"86",  -- 134
        16861 => X"96",  -- 150
        16862 => X"9D",  -- 157
        16863 => X"A0",  -- 160
        16864 => X"9B",  -- 155
        16865 => X"9B",  -- 155
        16866 => X"9B",  -- 155
        16867 => X"9C",  -- 156
        16868 => X"9D",  -- 157
        16869 => X"9D",  -- 157
        16870 => X"9A",  -- 154
        16871 => X"97",  -- 151
        16872 => X"93",  -- 147
        16873 => X"8C",  -- 140
        16874 => X"86",  -- 134
        16875 => X"83",  -- 131
        16876 => X"82",  -- 130
        16877 => X"80",  -- 128
        16878 => X"7C",  -- 124
        16879 => X"78",  -- 120
        16880 => X"72",  -- 114
        16881 => X"7B",  -- 123
        16882 => X"7C",  -- 124
        16883 => X"78",  -- 120
        16884 => X"6E",  -- 110
        16885 => X"5C",  -- 92
        16886 => X"56",  -- 86
        16887 => X"62",  -- 98
        16888 => X"68",  -- 104
        16889 => X"76",  -- 118
        16890 => X"82",  -- 130
        16891 => X"8A",  -- 138
        16892 => X"8F",  -- 143
        16893 => X"96",  -- 150
        16894 => X"9A",  -- 154
        16895 => X"9D",  -- 157
        16896 => X"9D",  -- 157
        16897 => X"9E",  -- 158
        16898 => X"A0",  -- 160
        16899 => X"A4",  -- 164
        16900 => X"AC",  -- 172
        16901 => X"AE",  -- 174
        16902 => X"AB",  -- 171
        16903 => X"A5",  -- 165
        16904 => X"A6",  -- 166
        16905 => X"9F",  -- 159
        16906 => X"95",  -- 149
        16907 => X"8B",  -- 139
        16908 => X"84",  -- 132
        16909 => X"80",  -- 128
        16910 => X"7C",  -- 124
        16911 => X"7A",  -- 122
        16912 => X"79",  -- 121
        16913 => X"7C",  -- 124
        16914 => X"7F",  -- 127
        16915 => X"7E",  -- 126
        16916 => X"74",  -- 116
        16917 => X"5E",  -- 94
        16918 => X"43",  -- 67
        16919 => X"2F",  -- 47
        16920 => X"23",  -- 35
        16921 => X"28",  -- 40
        16922 => X"3E",  -- 62
        16923 => X"5F",  -- 95
        16924 => X"72",  -- 114
        16925 => X"7B",  -- 123
        16926 => X"86",  -- 134
        16927 => X"94",  -- 148
        16928 => X"96",  -- 150
        16929 => X"97",  -- 151
        16930 => X"97",  -- 151
        16931 => X"9B",  -- 155
        16932 => X"A0",  -- 160
        16933 => X"9D",  -- 157
        16934 => X"86",  -- 134
        16935 => X"6C",  -- 108
        16936 => X"64",  -- 100
        16937 => X"70",  -- 112
        16938 => X"86",  -- 134
        16939 => X"9A",  -- 154
        16940 => X"A3",  -- 163
        16941 => X"A5",  -- 165
        16942 => X"AB",  -- 171
        16943 => X"B4",  -- 180
        16944 => X"B6",  -- 182
        16945 => X"B7",  -- 183
        16946 => X"B6",  -- 182
        16947 => X"B0",  -- 176
        16948 => X"B1",  -- 177
        16949 => X"B7",  -- 183
        16950 => X"BE",  -- 190
        16951 => X"C1",  -- 193
        16952 => X"BC",  -- 188
        16953 => X"B5",  -- 181
        16954 => X"B4",  -- 180
        16955 => X"BB",  -- 187
        16956 => X"BD",  -- 189
        16957 => X"B7",  -- 183
        16958 => X"B9",  -- 185
        16959 => X"C1",  -- 193
        16960 => X"7C",  -- 124
        16961 => X"7D",  -- 125
        16962 => X"7E",  -- 126
        16963 => X"7E",  -- 126
        16964 => X"7C",  -- 124
        16965 => X"7A",  -- 122
        16966 => X"77",  -- 119
        16967 => X"76",  -- 118
        16968 => X"75",  -- 117
        16969 => X"77",  -- 119
        16970 => X"77",  -- 119
        16971 => X"75",  -- 117
        16972 => X"73",  -- 115
        16973 => X"77",  -- 119
        16974 => X"7D",  -- 125
        16975 => X"85",  -- 133
        16976 => X"8C",  -- 140
        16977 => X"7C",  -- 124
        16978 => X"2C",  -- 44
        16979 => X"25",  -- 37
        16980 => X"42",  -- 66
        16981 => X"57",  -- 87
        16982 => X"54",  -- 84
        16983 => X"4A",  -- 74
        16984 => X"4A",  -- 74
        16985 => X"44",  -- 68
        16986 => X"40",  -- 64
        16987 => X"43",  -- 67
        16988 => X"44",  -- 68
        16989 => X"40",  -- 64
        16990 => X"3F",  -- 63
        16991 => X"42",  -- 66
        16992 => X"62",  -- 98
        16993 => X"6F",  -- 111
        16994 => X"6B",  -- 107
        16995 => X"58",  -- 88
        16996 => X"59",  -- 89
        16997 => X"6D",  -- 109
        16998 => X"72",  -- 114
        16999 => X"65",  -- 101
        17000 => X"56",  -- 86
        17001 => X"64",  -- 100
        17002 => X"5E",  -- 94
        17003 => X"4F",  -- 79
        17004 => X"4E",  -- 78
        17005 => X"53",  -- 83
        17006 => X"4E",  -- 78
        17007 => X"49",  -- 73
        17008 => X"4C",  -- 76
        17009 => X"57",  -- 87
        17010 => X"6B",  -- 107
        17011 => X"7A",  -- 122
        17012 => X"7B",  -- 123
        17013 => X"70",  -- 112
        17014 => X"65",  -- 101
        17015 => X"5F",  -- 95
        17016 => X"65",  -- 101
        17017 => X"84",  -- 132
        17018 => X"86",  -- 134
        17019 => X"81",  -- 129
        17020 => X"8F",  -- 143
        17021 => X"85",  -- 133
        17022 => X"5C",  -- 92
        17023 => X"40",  -- 64
        17024 => X"60",  -- 96
        17025 => X"71",  -- 113
        17026 => X"7F",  -- 127
        17027 => X"7C",  -- 124
        17028 => X"6E",  -- 110
        17029 => X"44",  -- 68
        17030 => X"18",  -- 24
        17031 => X"1E",  -- 30
        17032 => X"0C",  -- 12
        17033 => X"05",  -- 5
        17034 => X"08",  -- 8
        17035 => X"09",  -- 9
        17036 => X"0D",  -- 13
        17037 => X"02",  -- 2
        17038 => X"0C",  -- 12
        17039 => X"18",  -- 24
        17040 => X"10",  -- 16
        17041 => X"0F",  -- 15
        17042 => X"10",  -- 16
        17043 => X"25",  -- 37
        17044 => X"18",  -- 24
        17045 => X"16",  -- 22
        17046 => X"1B",  -- 27
        17047 => X"36",  -- 54
        17048 => X"41",  -- 65
        17049 => X"2F",  -- 47
        17050 => X"1A",  -- 26
        17051 => X"26",  -- 38
        17052 => X"3C",  -- 60
        17053 => X"2F",  -- 47
        17054 => X"2C",  -- 44
        17055 => X"50",  -- 80
        17056 => X"47",  -- 71
        17057 => X"4E",  -- 78
        17058 => X"60",  -- 96
        17059 => X"55",  -- 85
        17060 => X"57",  -- 87
        17061 => X"77",  -- 119
        17062 => X"79",  -- 121
        17063 => X"61",  -- 97
        17064 => X"3C",  -- 60
        17065 => X"27",  -- 39
        17066 => X"31",  -- 49
        17067 => X"2F",  -- 47
        17068 => X"38",  -- 56
        17069 => X"34",  -- 52
        17070 => X"29",  -- 41
        17071 => X"19",  -- 25
        17072 => X"17",  -- 23
        17073 => X"1A",  -- 26
        17074 => X"17",  -- 23
        17075 => X"18",  -- 24
        17076 => X"1D",  -- 29
        17077 => X"18",  -- 24
        17078 => X"13",  -- 19
        17079 => X"19",  -- 25
        17080 => X"24",  -- 36
        17081 => X"21",  -- 33
        17082 => X"19",  -- 25
        17083 => X"26",  -- 38
        17084 => X"4F",  -- 79
        17085 => X"72",  -- 114
        17086 => X"7D",  -- 125
        17087 => X"7E",  -- 126
        17088 => X"54",  -- 84
        17089 => X"3A",  -- 58
        17090 => X"5B",  -- 91
        17091 => X"6B",  -- 107
        17092 => X"79",  -- 121
        17093 => X"67",  -- 103
        17094 => X"59",  -- 89
        17095 => X"47",  -- 71
        17096 => X"4C",  -- 76
        17097 => X"50",  -- 80
        17098 => X"53",  -- 83
        17099 => X"4A",  -- 74
        17100 => X"39",  -- 57
        17101 => X"35",  -- 53
        17102 => X"32",  -- 50
        17103 => X"2B",  -- 43
        17104 => X"3E",  -- 62
        17105 => X"3B",  -- 59
        17106 => X"4F",  -- 79
        17107 => X"58",  -- 88
        17108 => X"56",  -- 86
        17109 => X"69",  -- 105
        17110 => X"77",  -- 119
        17111 => X"63",  -- 99
        17112 => X"72",  -- 114
        17113 => X"5A",  -- 90
        17114 => X"60",  -- 96
        17115 => X"73",  -- 115
        17116 => X"6C",  -- 108
        17117 => X"59",  -- 89
        17118 => X"6B",  -- 107
        17119 => X"8F",  -- 143
        17120 => X"49",  -- 73
        17121 => X"67",  -- 103
        17122 => X"71",  -- 113
        17123 => X"5C",  -- 92
        17124 => X"4D",  -- 77
        17125 => X"48",  -- 72
        17126 => X"50",  -- 80
        17127 => X"59",  -- 89
        17128 => X"5A",  -- 90
        17129 => X"65",  -- 101
        17130 => X"64",  -- 100
        17131 => X"5F",  -- 95
        17132 => X"3D",  -- 61
        17133 => X"24",  -- 36
        17134 => X"9A",  -- 154
        17135 => X"AF",  -- 175
        17136 => X"98",  -- 152
        17137 => X"83",  -- 131
        17138 => X"71",  -- 113
        17139 => X"6C",  -- 108
        17140 => X"6E",  -- 110
        17141 => X"6F",  -- 111
        17142 => X"71",  -- 113
        17143 => X"75",  -- 117
        17144 => X"71",  -- 113
        17145 => X"67",  -- 103
        17146 => X"5F",  -- 95
        17147 => X"62",  -- 98
        17148 => X"6E",  -- 110
        17149 => X"78",  -- 120
        17150 => X"78",  -- 120
        17151 => X"75",  -- 117
        17152 => X"7D",  -- 125
        17153 => X"7C",  -- 124
        17154 => X"7C",  -- 124
        17155 => X"7C",  -- 124
        17156 => X"7D",  -- 125
        17157 => X"81",  -- 129
        17158 => X"83",  -- 131
        17159 => X"85",  -- 133
        17160 => X"76",  -- 118
        17161 => X"77",  -- 119
        17162 => X"79",  -- 121
        17163 => X"78",  -- 120
        17164 => X"7D",  -- 125
        17165 => X"85",  -- 133
        17166 => X"89",  -- 137
        17167 => X"88",  -- 136
        17168 => X"98",  -- 152
        17169 => X"97",  -- 151
        17170 => X"98",  -- 152
        17171 => X"9A",  -- 154
        17172 => X"99",  -- 153
        17173 => X"95",  -- 149
        17174 => X"92",  -- 146
        17175 => X"93",  -- 147
        17176 => X"8D",  -- 141
        17177 => X"83",  -- 131
        17178 => X"79",  -- 121
        17179 => X"7B",  -- 123
        17180 => X"87",  -- 135
        17181 => X"96",  -- 150
        17182 => X"9E",  -- 158
        17183 => X"A3",  -- 163
        17184 => X"98",  -- 152
        17185 => X"9B",  -- 155
        17186 => X"9F",  -- 159
        17187 => X"9F",  -- 159
        17188 => X"A1",  -- 161
        17189 => X"9E",  -- 158
        17190 => X"9A",  -- 154
        17191 => X"92",  -- 146
        17192 => X"95",  -- 149
        17193 => X"8F",  -- 143
        17194 => X"8A",  -- 138
        17195 => X"88",  -- 136
        17196 => X"85",  -- 133
        17197 => X"80",  -- 128
        17198 => X"7B",  -- 123
        17199 => X"7A",  -- 122
        17200 => X"7A",  -- 122
        17201 => X"7C",  -- 124
        17202 => X"78",  -- 120
        17203 => X"75",  -- 117
        17204 => X"72",  -- 114
        17205 => X"61",  -- 97
        17206 => X"51",  -- 81
        17207 => X"51",  -- 81
        17208 => X"5F",  -- 95
        17209 => X"71",  -- 113
        17210 => X"85",  -- 133
        17211 => X"8D",  -- 141
        17212 => X"93",  -- 147
        17213 => X"99",  -- 153
        17214 => X"9C",  -- 156
        17215 => X"9B",  -- 155
        17216 => X"9C",  -- 156
        17217 => X"9E",  -- 158
        17218 => X"A2",  -- 162
        17219 => X"A6",  -- 166
        17220 => X"AB",  -- 171
        17221 => X"AB",  -- 171
        17222 => X"A7",  -- 167
        17223 => X"A3",  -- 163
        17224 => X"9E",  -- 158
        17225 => X"9A",  -- 154
        17226 => X"96",  -- 150
        17227 => X"8F",  -- 143
        17228 => X"87",  -- 135
        17229 => X"80",  -- 128
        17230 => X"7C",  -- 124
        17231 => X"7A",  -- 122
        17232 => X"82",  -- 130
        17233 => X"7F",  -- 127
        17234 => X"7F",  -- 127
        17235 => X"7F",  -- 127
        17236 => X"75",  -- 117
        17237 => X"5A",  -- 90
        17238 => X"38",  -- 56
        17239 => X"20",  -- 32
        17240 => X"18",  -- 24
        17241 => X"25",  -- 37
        17242 => X"44",  -- 68
        17243 => X"67",  -- 103
        17244 => X"7A",  -- 122
        17245 => X"80",  -- 128
        17246 => X"89",  -- 137
        17247 => X"94",  -- 148
        17248 => X"8E",  -- 142
        17249 => X"92",  -- 146
        17250 => X"94",  -- 148
        17251 => X"97",  -- 151
        17252 => X"9A",  -- 154
        17253 => X"91",  -- 145
        17254 => X"72",  -- 114
        17255 => X"55",  -- 85
        17256 => X"57",  -- 87
        17257 => X"6D",  -- 109
        17258 => X"88",  -- 136
        17259 => X"99",  -- 153
        17260 => X"A1",  -- 161
        17261 => X"A6",  -- 166
        17262 => X"AA",  -- 170
        17263 => X"AC",  -- 172
        17264 => X"B1",  -- 177
        17265 => X"B5",  -- 181
        17266 => X"B4",  -- 180
        17267 => X"AD",  -- 173
        17268 => X"AF",  -- 175
        17269 => X"B7",  -- 183
        17270 => X"BD",  -- 189
        17271 => X"BD",  -- 189
        17272 => X"B8",  -- 184
        17273 => X"B2",  -- 178
        17274 => X"B3",  -- 179
        17275 => X"BB",  -- 187
        17276 => X"BC",  -- 188
        17277 => X"B6",  -- 182
        17278 => X"BA",  -- 186
        17279 => X"C6",  -- 198
        17280 => X"81",  -- 129
        17281 => X"81",  -- 129
        17282 => X"80",  -- 128
        17283 => X"7F",  -- 127
        17284 => X"7D",  -- 125
        17285 => X"7D",  -- 125
        17286 => X"7D",  -- 125
        17287 => X"7D",  -- 125
        17288 => X"78",  -- 120
        17289 => X"7A",  -- 122
        17290 => X"7B",  -- 123
        17291 => X"7B",  -- 123
        17292 => X"7C",  -- 124
        17293 => X"7D",  -- 125
        17294 => X"80",  -- 128
        17295 => X"82",  -- 130
        17296 => X"8F",  -- 143
        17297 => X"69",  -- 105
        17298 => X"19",  -- 25
        17299 => X"28",  -- 40
        17300 => X"4F",  -- 79
        17301 => X"5A",  -- 90
        17302 => X"53",  -- 83
        17303 => X"55",  -- 85
        17304 => X"51",  -- 81
        17305 => X"49",  -- 73
        17306 => X"3F",  -- 63
        17307 => X"3C",  -- 60
        17308 => X"3F",  -- 63
        17309 => X"44",  -- 68
        17310 => X"4B",  -- 75
        17311 => X"4F",  -- 79
        17312 => X"59",  -- 89
        17313 => X"5A",  -- 90
        17314 => X"53",  -- 83
        17315 => X"51",  -- 81
        17316 => X"66",  -- 102
        17317 => X"7E",  -- 126
        17318 => X"7C",  -- 124
        17319 => X"6A",  -- 106
        17320 => X"5D",  -- 93
        17321 => X"6F",  -- 111
        17322 => X"6C",  -- 108
        17323 => X"58",  -- 88
        17324 => X"57",  -- 87
        17325 => X"5E",  -- 94
        17326 => X"51",  -- 81
        17327 => X"41",  -- 65
        17328 => X"53",  -- 83
        17329 => X"54",  -- 84
        17330 => X"57",  -- 87
        17331 => X"60",  -- 96
        17332 => X"72",  -- 114
        17333 => X"85",  -- 133
        17334 => X"90",  -- 144
        17335 => X"92",  -- 146
        17336 => X"64",  -- 100
        17337 => X"67",  -- 103
        17338 => X"73",  -- 115
        17339 => X"7C",  -- 124
        17340 => X"7C",  -- 124
        17341 => X"86",  -- 134
        17342 => X"7D",  -- 125
        17343 => X"60",  -- 96
        17344 => X"5D",  -- 93
        17345 => X"50",  -- 80
        17346 => X"6A",  -- 106
        17347 => X"69",  -- 105
        17348 => X"41",  -- 65
        17349 => X"20",  -- 32
        17350 => X"0C",  -- 12
        17351 => X"10",  -- 16
        17352 => X"10",  -- 16
        17353 => X"0A",  -- 10
        17354 => X"16",  -- 22
        17355 => X"13",  -- 19
        17356 => X"18",  -- 24
        17357 => X"09",  -- 9
        17358 => X"1D",  -- 29
        17359 => X"31",  -- 49
        17360 => X"36",  -- 54
        17361 => X"38",  -- 56
        17362 => X"35",  -- 53
        17363 => X"3E",  -- 62
        17364 => X"2E",  -- 46
        17365 => X"32",  -- 50
        17366 => X"45",  -- 69
        17367 => X"6B",  -- 107
        17368 => X"81",  -- 129
        17369 => X"6F",  -- 111
        17370 => X"57",  -- 87
        17371 => X"64",  -- 100
        17372 => X"76",  -- 118
        17373 => X"51",  -- 81
        17374 => X"2E",  -- 46
        17375 => X"3E",  -- 62
        17376 => X"3A",  -- 58
        17377 => X"31",  -- 49
        17378 => X"40",  -- 64
        17379 => X"4A",  -- 74
        17380 => X"4F",  -- 79
        17381 => X"56",  -- 86
        17382 => X"61",  -- 97
        17383 => X"7C",  -- 124
        17384 => X"6A",  -- 106
        17385 => X"56",  -- 86
        17386 => X"69",  -- 105
        17387 => X"66",  -- 102
        17388 => X"71",  -- 113
        17389 => X"6E",  -- 110
        17390 => X"5E",  -- 94
        17391 => X"40",  -- 64
        17392 => X"35",  -- 53
        17393 => X"33",  -- 51
        17394 => X"23",  -- 35
        17395 => X"19",  -- 25
        17396 => X"24",  -- 36
        17397 => X"22",  -- 34
        17398 => X"16",  -- 22
        17399 => X"16",  -- 22
        17400 => X"21",  -- 33
        17401 => X"28",  -- 40
        17402 => X"1B",  -- 27
        17403 => X"11",  -- 17
        17404 => X"27",  -- 39
        17405 => X"4D",  -- 77
        17406 => X"6C",  -- 108
        17407 => X"7C",  -- 124
        17408 => X"6A",  -- 106
        17409 => X"56",  -- 86
        17410 => X"6C",  -- 108
        17411 => X"73",  -- 115
        17412 => X"64",  -- 100
        17413 => X"5C",  -- 92
        17414 => X"56",  -- 86
        17415 => X"50",  -- 80
        17416 => X"59",  -- 89
        17417 => X"4B",  -- 75
        17418 => X"3A",  -- 58
        17419 => X"35",  -- 53
        17420 => X"36",  -- 54
        17421 => X"31",  -- 49
        17422 => X"32",  -- 50
        17423 => X"3C",  -- 60
        17424 => X"3F",  -- 63
        17425 => X"39",  -- 57
        17426 => X"58",  -- 88
        17427 => X"74",  -- 116
        17428 => X"74",  -- 116
        17429 => X"7C",  -- 124
        17430 => X"73",  -- 115
        17431 => X"4D",  -- 77
        17432 => X"7C",  -- 124
        17433 => X"69",  -- 105
        17434 => X"66",  -- 102
        17435 => X"5E",  -- 94
        17436 => X"69",  -- 105
        17437 => X"4E",  -- 78
        17438 => X"65",  -- 101
        17439 => X"7D",  -- 125
        17440 => X"6C",  -- 108
        17441 => X"67",  -- 103
        17442 => X"74",  -- 116
        17443 => X"5E",  -- 94
        17444 => X"51",  -- 81
        17445 => X"38",  -- 56
        17446 => X"4A",  -- 74
        17447 => X"53",  -- 83
        17448 => X"5B",  -- 91
        17449 => X"64",  -- 100
        17450 => X"67",  -- 103
        17451 => X"64",  -- 100
        17452 => X"5B",  -- 91
        17453 => X"28",  -- 40
        17454 => X"6A",  -- 106
        17455 => X"AF",  -- 175
        17456 => X"91",  -- 145
        17457 => X"7D",  -- 125
        17458 => X"6F",  -- 111
        17459 => X"71",  -- 113
        17460 => X"77",  -- 119
        17461 => X"77",  -- 119
        17462 => X"75",  -- 117
        17463 => X"74",  -- 116
        17464 => X"70",  -- 112
        17465 => X"69",  -- 105
        17466 => X"63",  -- 99
        17467 => X"68",  -- 104
        17468 => X"72",  -- 114
        17469 => X"77",  -- 119
        17470 => X"74",  -- 116
        17471 => X"6D",  -- 109
        17472 => X"72",  -- 114
        17473 => X"71",  -- 113
        17474 => X"72",  -- 114
        17475 => X"75",  -- 117
        17476 => X"7B",  -- 123
        17477 => X"80",  -- 128
        17478 => X"82",  -- 130
        17479 => X"82",  -- 130
        17480 => X"6D",  -- 109
        17481 => X"76",  -- 118
        17482 => X"7F",  -- 127
        17483 => X"85",  -- 133
        17484 => X"8A",  -- 138
        17485 => X"8F",  -- 143
        17486 => X"90",  -- 144
        17487 => X"8E",  -- 142
        17488 => X"94",  -- 148
        17489 => X"93",  -- 147
        17490 => X"97",  -- 151
        17491 => X"9A",  -- 154
        17492 => X"98",  -- 152
        17493 => X"90",  -- 144
        17494 => X"8C",  -- 140
        17495 => X"8C",  -- 140
        17496 => X"91",  -- 145
        17497 => X"8E",  -- 142
        17498 => X"89",  -- 137
        17499 => X"82",  -- 130
        17500 => X"7F",  -- 127
        17501 => X"86",  -- 134
        17502 => X"95",  -- 149
        17503 => X"A1",  -- 161
        17504 => X"9E",  -- 158
        17505 => X"A0",  -- 160
        17506 => X"9F",  -- 159
        17507 => X"9C",  -- 156
        17508 => X"9C",  -- 156
        17509 => X"9E",  -- 158
        17510 => X"9A",  -- 154
        17511 => X"95",  -- 149
        17512 => X"98",  -- 152
        17513 => X"93",  -- 147
        17514 => X"8F",  -- 143
        17515 => X"8C",  -- 140
        17516 => X"87",  -- 135
        17517 => X"7E",  -- 126
        17518 => X"79",  -- 121
        17519 => X"7A",  -- 122
        17520 => X"7C",  -- 124
        17521 => X"7D",  -- 125
        17522 => X"78",  -- 120
        17523 => X"76",  -- 118
        17524 => X"74",  -- 116
        17525 => X"64",  -- 100
        17526 => X"4F",  -- 79
        17527 => X"4A",  -- 74
        17528 => X"53",  -- 83
        17529 => X"67",  -- 103
        17530 => X"78",  -- 120
        17531 => X"7F",  -- 127
        17532 => X"85",  -- 133
        17533 => X"8C",  -- 140
        17534 => X"90",  -- 144
        17535 => X"8D",  -- 141
        17536 => X"96",  -- 150
        17537 => X"9A",  -- 154
        17538 => X"A1",  -- 161
        17539 => X"A7",  -- 167
        17540 => X"A9",  -- 169
        17541 => X"A7",  -- 167
        17542 => X"A4",  -- 164
        17543 => X"A1",  -- 161
        17544 => X"9F",  -- 159
        17545 => X"9E",  -- 158
        17546 => X"9C",  -- 156
        17547 => X"96",  -- 150
        17548 => X"8E",  -- 142
        17549 => X"88",  -- 136
        17550 => X"84",  -- 132
        17551 => X"84",  -- 132
        17552 => X"86",  -- 134
        17553 => X"81",  -- 129
        17554 => X"80",  -- 128
        17555 => X"81",  -- 129
        17556 => X"73",  -- 115
        17557 => X"51",  -- 81
        17558 => X"2E",  -- 46
        17559 => X"1B",  -- 27
        17560 => X"18",  -- 24
        17561 => X"29",  -- 41
        17562 => X"47",  -- 71
        17563 => X"65",  -- 101
        17564 => X"78",  -- 120
        17565 => X"80",  -- 128
        17566 => X"86",  -- 134
        17567 => X"8B",  -- 139
        17568 => X"88",  -- 136
        17569 => X"8D",  -- 141
        17570 => X"90",  -- 144
        17571 => X"8F",  -- 143
        17572 => X"8E",  -- 142
        17573 => X"85",  -- 133
        17574 => X"6B",  -- 107
        17575 => X"54",  -- 84
        17576 => X"59",  -- 89
        17577 => X"75",  -- 117
        17578 => X"90",  -- 144
        17579 => X"9A",  -- 154
        17580 => X"A0",  -- 160
        17581 => X"AA",  -- 170
        17582 => X"AC",  -- 172
        17583 => X"A7",  -- 167
        17584 => X"AE",  -- 174
        17585 => X"B2",  -- 178
        17586 => X"B2",  -- 178
        17587 => X"AB",  -- 171
        17588 => X"AC",  -- 172
        17589 => X"B5",  -- 181
        17590 => X"B9",  -- 185
        17591 => X"B7",  -- 183
        17592 => X"B6",  -- 182
        17593 => X"B3",  -- 179
        17594 => X"B7",  -- 183
        17595 => X"BE",  -- 190
        17596 => X"BC",  -- 188
        17597 => X"B6",  -- 182
        17598 => X"B9",  -- 185
        17599 => X"C5",  -- 197
        17600 => X"87",  -- 135
        17601 => X"85",  -- 133
        17602 => X"81",  -- 129
        17603 => X"7D",  -- 125
        17604 => X"7B",  -- 123
        17605 => X"7C",  -- 124
        17606 => X"7D",  -- 125
        17607 => X"7C",  -- 124
        17608 => X"78",  -- 120
        17609 => X"7B",  -- 123
        17610 => X"7D",  -- 125
        17611 => X"81",  -- 129
        17612 => X"82",  -- 130
        17613 => X"83",  -- 131
        17614 => X"82",  -- 130
        17615 => X"82",  -- 130
        17616 => X"81",  -- 129
        17617 => X"87",  -- 135
        17618 => X"4F",  -- 79
        17619 => X"4C",  -- 76
        17620 => X"56",  -- 86
        17621 => X"59",  -- 89
        17622 => X"5E",  -- 94
        17623 => X"64",  -- 100
        17624 => X"56",  -- 86
        17625 => X"4D",  -- 77
        17626 => X"3E",  -- 62
        17627 => X"36",  -- 54
        17628 => X"38",  -- 56
        17629 => X"45",  -- 69
        17630 => X"50",  -- 80
        17631 => X"54",  -- 84
        17632 => X"5C",  -- 92
        17633 => X"51",  -- 81
        17634 => X"5A",  -- 90
        17635 => X"75",  -- 117
        17636 => X"82",  -- 130
        17637 => X"6D",  -- 109
        17638 => X"4D",  -- 77
        17639 => X"39",  -- 57
        17640 => X"48",  -- 72
        17641 => X"6C",  -- 108
        17642 => X"75",  -- 117
        17643 => X"67",  -- 103
        17644 => X"65",  -- 101
        17645 => X"6E",  -- 110
        17646 => X"64",  -- 100
        17647 => X"52",  -- 82
        17648 => X"34",  -- 52
        17649 => X"3C",  -- 60
        17650 => X"43",  -- 67
        17651 => X"4B",  -- 75
        17652 => X"5D",  -- 93
        17653 => X"75",  -- 117
        17654 => X"89",  -- 137
        17655 => X"90",  -- 144
        17656 => X"8E",  -- 142
        17657 => X"5A",  -- 90
        17658 => X"64",  -- 100
        17659 => X"7C",  -- 124
        17660 => X"68",  -- 104
        17661 => X"76",  -- 118
        17662 => X"98",  -- 152
        17663 => X"8C",  -- 140
        17664 => X"8C",  -- 140
        17665 => X"54",  -- 84
        17666 => X"68",  -- 104
        17667 => X"64",  -- 100
        17668 => X"28",  -- 40
        17669 => X"14",  -- 20
        17670 => X"14",  -- 20
        17671 => X"0E",  -- 14
        17672 => X"0F",  -- 15
        17673 => X"09",  -- 9
        17674 => X"16",  -- 22
        17675 => X"19",  -- 25
        17676 => X"2F",  -- 47
        17677 => X"32",  -- 50
        17678 => X"53",  -- 83
        17679 => X"68",  -- 104
        17680 => X"69",  -- 105
        17681 => X"72",  -- 114
        17682 => X"73",  -- 115
        17683 => X"7A",  -- 122
        17684 => X"6B",  -- 107
        17685 => X"71",  -- 113
        17686 => X"7C",  -- 124
        17687 => X"93",  -- 147
        17688 => X"96",  -- 150
        17689 => X"93",  -- 147
        17690 => X"75",  -- 117
        17691 => X"6C",  -- 108
        17692 => X"7E",  -- 126
        17693 => X"65",  -- 101
        17694 => X"35",  -- 53
        17695 => X"2E",  -- 46
        17696 => X"2A",  -- 42
        17697 => X"23",  -- 35
        17698 => X"24",  -- 36
        17699 => X"1B",  -- 27
        17700 => X"1A",  -- 26
        17701 => X"20",  -- 32
        17702 => X"38",  -- 56
        17703 => X"6A",  -- 106
        17704 => X"81",  -- 129
        17705 => X"71",  -- 113
        17706 => X"84",  -- 132
        17707 => X"78",  -- 120
        17708 => X"80",  -- 128
        17709 => X"82",  -- 130
        17710 => X"81",  -- 129
        17711 => X"6C",  -- 108
        17712 => X"6A",  -- 106
        17713 => X"62",  -- 98
        17714 => X"44",  -- 68
        17715 => X"30",  -- 48
        17716 => X"39",  -- 57
        17717 => X"39",  -- 57
        17718 => X"27",  -- 39
        17719 => X"21",  -- 33
        17720 => X"22",  -- 34
        17721 => X"1A",  -- 26
        17722 => X"13",  -- 19
        17723 => X"16",  -- 22
        17724 => X"1C",  -- 28
        17725 => X"27",  -- 39
        17726 => X"53",  -- 83
        17727 => X"8B",  -- 139
        17728 => X"86",  -- 134
        17729 => X"75",  -- 117
        17730 => X"79",  -- 121
        17731 => X"78",  -- 120
        17732 => X"55",  -- 85
        17733 => X"5E",  -- 94
        17734 => X"59",  -- 89
        17735 => X"57",  -- 87
        17736 => X"4D",  -- 77
        17737 => X"41",  -- 65
        17738 => X"32",  -- 50
        17739 => X"34",  -- 52
        17740 => X"39",  -- 57
        17741 => X"2C",  -- 44
        17742 => X"36",  -- 54
        17743 => X"5B",  -- 91
        17744 => X"6B",  -- 107
        17745 => X"58",  -- 88
        17746 => X"63",  -- 99
        17747 => X"68",  -- 104
        17748 => X"5A",  -- 90
        17749 => X"69",  -- 105
        17750 => X"81",  -- 129
        17751 => X"75",  -- 117
        17752 => X"47",  -- 71
        17753 => X"7B",  -- 123
        17754 => X"76",  -- 118
        17755 => X"6E",  -- 110
        17756 => X"84",  -- 132
        17757 => X"5C",  -- 92
        17758 => X"84",  -- 132
        17759 => X"65",  -- 101
        17760 => X"65",  -- 101
        17761 => X"50",  -- 80
        17762 => X"5B",  -- 91
        17763 => X"42",  -- 66
        17764 => X"46",  -- 70
        17765 => X"37",  -- 55
        17766 => X"5C",  -- 92
        17767 => X"5F",  -- 95
        17768 => X"6F",  -- 111
        17769 => X"67",  -- 103
        17770 => X"6A",  -- 106
        17771 => X"66",  -- 102
        17772 => X"72",  -- 114
        17773 => X"39",  -- 57
        17774 => X"44",  -- 68
        17775 => X"A1",  -- 161
        17776 => X"9E",  -- 158
        17777 => X"8A",  -- 138
        17778 => X"77",  -- 119
        17779 => X"6E",  -- 110
        17780 => X"6B",  -- 107
        17781 => X"67",  -- 103
        17782 => X"6D",  -- 109
        17783 => X"75",  -- 117
        17784 => X"70",  -- 112
        17785 => X"72",  -- 114
        17786 => X"74",  -- 116
        17787 => X"73",  -- 115
        17788 => X"71",  -- 113
        17789 => X"72",  -- 114
        17790 => X"73",  -- 115
        17791 => X"75",  -- 117
        17792 => X"69",  -- 105
        17793 => X"69",  -- 105
        17794 => X"6D",  -- 109
        17795 => X"76",  -- 118
        17796 => X"80",  -- 128
        17797 => X"85",  -- 133
        17798 => X"83",  -- 131
        17799 => X"7F",  -- 127
        17800 => X"84",  -- 132
        17801 => X"89",  -- 137
        17802 => X"8D",  -- 141
        17803 => X"8D",  -- 141
        17804 => X"8E",  -- 142
        17805 => X"96",  -- 150
        17806 => X"9D",  -- 157
        17807 => X"A0",  -- 160
        17808 => X"9C",  -- 156
        17809 => X"9D",  -- 157
        17810 => X"A0",  -- 160
        17811 => X"A4",  -- 164
        17812 => X"A0",  -- 160
        17813 => X"95",  -- 149
        17814 => X"8E",  -- 142
        17815 => X"8F",  -- 143
        17816 => X"95",  -- 149
        17817 => X"96",  -- 150
        17818 => X"8E",  -- 142
        17819 => X"7B",  -- 123
        17820 => X"6A",  -- 106
        17821 => X"6E",  -- 110
        17822 => X"84",  -- 132
        17823 => X"98",  -- 152
        17824 => X"AA",  -- 170
        17825 => X"A6",  -- 166
        17826 => X"9F",  -- 159
        17827 => X"95",  -- 149
        17828 => X"93",  -- 147
        17829 => X"99",  -- 153
        17830 => X"9D",  -- 157
        17831 => X"9B",  -- 155
        17832 => X"97",  -- 151
        17833 => X"93",  -- 147
        17834 => X"90",  -- 144
        17835 => X"8D",  -- 141
        17836 => X"84",  -- 132
        17837 => X"79",  -- 121
        17838 => X"74",  -- 116
        17839 => X"76",  -- 118
        17840 => X"75",  -- 117
        17841 => X"7D",  -- 125
        17842 => X"7E",  -- 126
        17843 => X"7B",  -- 123
        17844 => X"74",  -- 116
        17845 => X"61",  -- 97
        17846 => X"50",  -- 80
        17847 => X"4D",  -- 77
        17848 => X"5B",  -- 91
        17849 => X"6C",  -- 108
        17850 => X"78",  -- 120
        17851 => X"79",  -- 121
        17852 => X"7D",  -- 125
        17853 => X"86",  -- 134
        17854 => X"8E",  -- 142
        17855 => X"8E",  -- 142
        17856 => X"91",  -- 145
        17857 => X"95",  -- 149
        17858 => X"9E",  -- 158
        17859 => X"A6",  -- 166
        17860 => X"A6",  -- 166
        17861 => X"A4",  -- 164
        17862 => X"A0",  -- 160
        17863 => X"9F",  -- 159
        17864 => X"A4",  -- 164
        17865 => X"A2",  -- 162
        17866 => X"9E",  -- 158
        17867 => X"95",  -- 149
        17868 => X"8D",  -- 141
        17869 => X"89",  -- 137
        17870 => X"89",  -- 137
        17871 => X"8A",  -- 138
        17872 => X"8B",  -- 139
        17873 => X"85",  -- 133
        17874 => X"85",  -- 133
        17875 => X"86",  -- 134
        17876 => X"76",  -- 118
        17877 => X"52",  -- 82
        17878 => X"32",  -- 50
        17879 => X"23",  -- 35
        17880 => X"27",  -- 39
        17881 => X"33",  -- 51
        17882 => X"4B",  -- 75
        17883 => X"64",  -- 100
        17884 => X"77",  -- 119
        17885 => X"81",  -- 129
        17886 => X"86",  -- 134
        17887 => X"88",  -- 136
        17888 => X"8C",  -- 140
        17889 => X"91",  -- 145
        17890 => X"93",  -- 147
        17891 => X"8E",  -- 142
        17892 => X"8C",  -- 140
        17893 => X"86",  -- 134
        17894 => X"79",  -- 121
        17895 => X"6B",  -- 107
        17896 => X"6C",  -- 108
        17897 => X"89",  -- 137
        17898 => X"9E",  -- 158
        17899 => X"9F",  -- 159
        17900 => X"A4",  -- 164
        17901 => X"B1",  -- 177
        17902 => X"B2",  -- 178
        17903 => X"AA",  -- 170
        17904 => X"AD",  -- 173
        17905 => X"B3",  -- 179
        17906 => X"B2",  -- 178
        17907 => X"AB",  -- 171
        17908 => X"AC",  -- 172
        17909 => X"B6",  -- 182
        17910 => X"BA",  -- 186
        17911 => X"B6",  -- 182
        17912 => X"B4",  -- 180
        17913 => X"B2",  -- 178
        17914 => X"B7",  -- 183
        17915 => X"BE",  -- 190
        17916 => X"BA",  -- 186
        17917 => X"B0",  -- 176
        17918 => X"B1",  -- 177
        17919 => X"BC",  -- 188
        17920 => X"8A",  -- 138
        17921 => X"8A",  -- 138
        17922 => X"88",  -- 136
        17923 => X"82",  -- 130
        17924 => X"7B",  -- 123
        17925 => X"78",  -- 120
        17926 => X"7B",  -- 123
        17927 => X"80",  -- 128
        17928 => X"7B",  -- 123
        17929 => X"7D",  -- 125
        17930 => X"82",  -- 130
        17931 => X"87",  -- 135
        17932 => X"8B",  -- 139
        17933 => X"8D",  -- 141
        17934 => X"8D",  -- 141
        17935 => X"8D",  -- 141
        17936 => X"8F",  -- 143
        17937 => X"8D",  -- 141
        17938 => X"68",  -- 104
        17939 => X"2A",  -- 42
        17940 => X"4D",  -- 77
        17941 => X"4F",  -- 79
        17942 => X"6B",  -- 107
        17943 => X"67",  -- 103
        17944 => X"57",  -- 87
        17945 => X"52",  -- 82
        17946 => X"45",  -- 69
        17947 => X"38",  -- 56
        17948 => X"3A",  -- 58
        17949 => X"4A",  -- 74
        17950 => X"52",  -- 82
        17951 => X"51",  -- 81
        17952 => X"67",  -- 103
        17953 => X"6E",  -- 110
        17954 => X"7B",  -- 123
        17955 => X"84",  -- 132
        17956 => X"84",  -- 132
        17957 => X"60",  -- 96
        17958 => X"4A",  -- 74
        17959 => X"50",  -- 80
        17960 => X"51",  -- 81
        17961 => X"46",  -- 70
        17962 => X"50",  -- 80
        17963 => X"64",  -- 100
        17964 => X"6A",  -- 106
        17965 => X"65",  -- 101
        17966 => X"61",  -- 97
        17967 => X"5F",  -- 95
        17968 => X"49",  -- 73
        17969 => X"53",  -- 83
        17970 => X"3D",  -- 61
        17971 => X"38",  -- 56
        17972 => X"4D",  -- 77
        17973 => X"5F",  -- 95
        17974 => X"6F",  -- 111
        17975 => X"79",  -- 121
        17976 => X"92",  -- 146
        17977 => X"8D",  -- 141
        17978 => X"65",  -- 101
        17979 => X"5D",  -- 93
        17980 => X"64",  -- 100
        17981 => X"71",  -- 113
        17982 => X"6D",  -- 109
        17983 => X"80",  -- 128
        17984 => X"85",  -- 133
        17985 => X"92",  -- 146
        17986 => X"70",  -- 112
        17987 => X"38",  -- 56
        17988 => X"27",  -- 39
        17989 => X"0D",  -- 13
        17990 => X"18",  -- 24
        17991 => X"0B",  -- 11
        17992 => X"1F",  -- 31
        17993 => X"2E",  -- 46
        17994 => X"4E",  -- 78
        17995 => X"46",  -- 70
        17996 => X"6B",  -- 107
        17997 => X"76",  -- 118
        17998 => X"91",  -- 145
        17999 => X"87",  -- 135
        18000 => X"88",  -- 136
        18001 => X"90",  -- 144
        18002 => X"8E",  -- 142
        18003 => X"83",  -- 131
        18004 => X"80",  -- 128
        18005 => X"83",  -- 131
        18006 => X"83",  -- 131
        18007 => X"7B",  -- 123
        18008 => X"68",  -- 104
        18009 => X"8A",  -- 138
        18010 => X"6C",  -- 108
        18011 => X"6C",  -- 108
        18012 => X"5E",  -- 94
        18013 => X"28",  -- 40
        18014 => X"23",  -- 35
        18015 => X"1D",  -- 29
        18016 => X"1D",  -- 29
        18017 => X"13",  -- 19
        18018 => X"0F",  -- 15
        18019 => X"1A",  -- 26
        18020 => X"0F",  -- 15
        18021 => X"10",  -- 16
        18022 => X"1B",  -- 27
        18023 => X"4C",  -- 76
        18024 => X"5D",  -- 93
        18025 => X"5B",  -- 91
        18026 => X"59",  -- 89
        18027 => X"5A",  -- 90
        18028 => X"68",  -- 104
        18029 => X"81",  -- 129
        18030 => X"88",  -- 136
        18031 => X"7C",  -- 124
        18032 => X"86",  -- 134
        18033 => X"8C",  -- 140
        18034 => X"82",  -- 130
        18035 => X"71",  -- 113
        18036 => X"69",  -- 105
        18037 => X"5D",  -- 93
        18038 => X"42",  -- 66
        18039 => X"2F",  -- 47
        18040 => X"25",  -- 37
        18041 => X"17",  -- 23
        18042 => X"10",  -- 16
        18043 => X"19",  -- 25
        18044 => X"1B",  -- 27
        18045 => X"18",  -- 24
        18046 => X"3A",  -- 58
        18047 => X"70",  -- 112
        18048 => X"8B",  -- 139
        18049 => X"78",  -- 120
        18050 => X"6E",  -- 110
        18051 => X"6B",  -- 107
        18052 => X"60",  -- 96
        18053 => X"58",  -- 88
        18054 => X"57",  -- 87
        18055 => X"54",  -- 84
        18056 => X"47",  -- 71
        18057 => X"31",  -- 49
        18058 => X"36",  -- 54
        18059 => X"30",  -- 48
        18060 => X"2F",  -- 47
        18061 => X"2C",  -- 44
        18062 => X"3E",  -- 62
        18063 => X"38",  -- 56
        18064 => X"5C",  -- 92
        18065 => X"57",  -- 87
        18066 => X"63",  -- 99
        18067 => X"6F",  -- 111
        18068 => X"64",  -- 100
        18069 => X"4D",  -- 77
        18070 => X"5D",  -- 93
        18071 => X"7F",  -- 127
        18072 => X"4E",  -- 78
        18073 => X"42",  -- 66
        18074 => X"94",  -- 148
        18075 => X"89",  -- 137
        18076 => X"87",  -- 135
        18077 => X"78",  -- 120
        18078 => X"8E",  -- 142
        18079 => X"66",  -- 102
        18080 => X"64",  -- 100
        18081 => X"37",  -- 55
        18082 => X"4E",  -- 78
        18083 => X"37",  -- 55
        18084 => X"4F",  -- 79
        18085 => X"51",  -- 81
        18086 => X"57",  -- 87
        18087 => X"66",  -- 102
        18088 => X"65",  -- 101
        18089 => X"5C",  -- 92
        18090 => X"65",  -- 101
        18091 => X"6A",  -- 106
        18092 => X"76",  -- 118
        18093 => X"57",  -- 87
        18094 => X"49",  -- 73
        18095 => X"A0",  -- 160
        18096 => X"A9",  -- 169
        18097 => X"8E",  -- 142
        18098 => X"76",  -- 118
        18099 => X"73",  -- 115
        18100 => X"7B",  -- 123
        18101 => X"7C",  -- 124
        18102 => X"7A",  -- 122
        18103 => X"79",  -- 121
        18104 => X"7E",  -- 126
        18105 => X"7E",  -- 126
        18106 => X"7F",  -- 127
        18107 => X"7D",  -- 125
        18108 => X"7B",  -- 123
        18109 => X"78",  -- 120
        18110 => X"76",  -- 118
        18111 => X"76",  -- 118
        18112 => X"68",  -- 104
        18113 => X"6B",  -- 107
        18114 => X"6D",  -- 109
        18115 => X"6D",  -- 109
        18116 => X"73",  -- 115
        18117 => X"7E",  -- 126
        18118 => X"85",  -- 133
        18119 => X"86",  -- 134
        18120 => X"88",  -- 136
        18121 => X"82",  -- 130
        18122 => X"81",  -- 129
        18123 => X"88",  -- 136
        18124 => X"96",  -- 150
        18125 => X"A2",  -- 162
        18126 => X"A4",  -- 164
        18127 => X"A2",  -- 162
        18128 => X"A2",  -- 162
        18129 => X"A8",  -- 168
        18130 => X"AE",  -- 174
        18131 => X"AC",  -- 172
        18132 => X"A3",  -- 163
        18133 => X"9D",  -- 157
        18134 => X"9D",  -- 157
        18135 => X"A1",  -- 161
        18136 => X"9F",  -- 159
        18137 => X"A8",  -- 168
        18138 => X"A0",  -- 160
        18139 => X"80",  -- 128
        18140 => X"6A",  -- 106
        18141 => X"70",  -- 112
        18142 => X"8B",  -- 139
        18143 => X"A0",  -- 160
        18144 => X"A8",  -- 168
        18145 => X"A1",  -- 161
        18146 => X"99",  -- 153
        18147 => X"98",  -- 152
        18148 => X"99",  -- 153
        18149 => X"9C",  -- 156
        18150 => X"9C",  -- 156
        18151 => X"9C",  -- 156
        18152 => X"97",  -- 151
        18153 => X"9A",  -- 154
        18154 => X"95",  -- 149
        18155 => X"89",  -- 137
        18156 => X"80",  -- 128
        18157 => X"7F",  -- 127
        18158 => X"7B",  -- 123
        18159 => X"75",  -- 117
        18160 => X"7A",  -- 122
        18161 => X"75",  -- 117
        18162 => X"79",  -- 121
        18163 => X"7E",  -- 126
        18164 => X"74",  -- 116
        18165 => X"60",  -- 96
        18166 => X"56",  -- 86
        18167 => X"59",  -- 89
        18168 => X"5F",  -- 95
        18169 => X"62",  -- 98
        18170 => X"68",  -- 104
        18171 => X"6F",  -- 111
        18172 => X"78",  -- 120
        18173 => X"80",  -- 128
        18174 => X"81",  -- 129
        18175 => X"83",  -- 131
        18176 => X"8A",  -- 138
        18177 => X"8D",  -- 141
        18178 => X"92",  -- 146
        18179 => X"9A",  -- 154
        18180 => X"A0",  -- 160
        18181 => X"A6",  -- 166
        18182 => X"A7",  -- 167
        18183 => X"A9",  -- 169
        18184 => X"A9",  -- 169
        18185 => X"A9",  -- 169
        18186 => X"A3",  -- 163
        18187 => X"98",  -- 152
        18188 => X"91",  -- 145
        18189 => X"92",  -- 146
        18190 => X"92",  -- 146
        18191 => X"90",  -- 144
        18192 => X"96",  -- 150
        18193 => X"8A",  -- 138
        18194 => X"89",  -- 137
        18195 => X"88",  -- 136
        18196 => X"6F",  -- 111
        18197 => X"42",  -- 66
        18198 => X"26",  -- 38
        18199 => X"21",  -- 33
        18200 => X"22",  -- 34
        18201 => X"30",  -- 48
        18202 => X"4B",  -- 75
        18203 => X"69",  -- 105
        18204 => X"7C",  -- 124
        18205 => X"86",  -- 134
        18206 => X"90",  -- 144
        18207 => X"99",  -- 153
        18208 => X"92",  -- 146
        18209 => X"94",  -- 148
        18210 => X"90",  -- 144
        18211 => X"90",  -- 144
        18212 => X"93",  -- 147
        18213 => X"83",  -- 131
        18214 => X"6D",  -- 109
        18215 => X"66",  -- 102
        18216 => X"76",  -- 118
        18217 => X"90",  -- 144
        18218 => X"A1",  -- 161
        18219 => X"A6",  -- 166
        18220 => X"AB",  -- 171
        18221 => X"AE",  -- 174
        18222 => X"AD",  -- 173
        18223 => X"B0",  -- 176
        18224 => X"B1",  -- 177
        18225 => X"B1",  -- 177
        18226 => X"AB",  -- 171
        18227 => X"A8",  -- 168
        18228 => X"B2",  -- 178
        18229 => X"BE",  -- 190
        18230 => X"BD",  -- 189
        18231 => X"B4",  -- 180
        18232 => X"B8",  -- 184
        18233 => X"BE",  -- 190
        18234 => X"BF",  -- 191
        18235 => X"C0",  -- 192
        18236 => X"BD",  -- 189
        18237 => X"B1",  -- 177
        18238 => X"A7",  -- 167
        18239 => X"AD",  -- 173
        18240 => X"88",  -- 136
        18241 => X"88",  -- 136
        18242 => X"85",  -- 133
        18243 => X"81",  -- 129
        18244 => X"7A",  -- 122
        18245 => X"79",  -- 121
        18246 => X"7A",  -- 122
        18247 => X"7E",  -- 126
        18248 => X"81",  -- 129
        18249 => X"84",  -- 132
        18250 => X"8A",  -- 138
        18251 => X"90",  -- 144
        18252 => X"94",  -- 148
        18253 => X"97",  -- 151
        18254 => X"97",  -- 151
        18255 => X"97",  -- 151
        18256 => X"8C",  -- 140
        18257 => X"7F",  -- 127
        18258 => X"2D",  -- 45
        18259 => X"3A",  -- 58
        18260 => X"49",  -- 73
        18261 => X"47",  -- 71
        18262 => X"4D",  -- 77
        18263 => X"5E",  -- 94
        18264 => X"57",  -- 87
        18265 => X"55",  -- 85
        18266 => X"4B",  -- 75
        18267 => X"3D",  -- 61
        18268 => X"3C",  -- 60
        18269 => X"4D",  -- 77
        18270 => X"5C",  -- 92
        18271 => X"63",  -- 99
        18272 => X"6D",  -- 109
        18273 => X"7A",  -- 122
        18274 => X"88",  -- 136
        18275 => X"90",  -- 144
        18276 => X"76",  -- 118
        18277 => X"6D",  -- 109
        18278 => X"55",  -- 85
        18279 => X"40",  -- 64
        18280 => X"2C",  -- 44
        18281 => X"3B",  -- 59
        18282 => X"5B",  -- 91
        18283 => X"74",  -- 116
        18284 => X"70",  -- 112
        18285 => X"61",  -- 97
        18286 => X"52",  -- 82
        18287 => X"49",  -- 73
        18288 => X"71",  -- 113
        18289 => X"7E",  -- 126
        18290 => X"66",  -- 102
        18291 => X"4C",  -- 76
        18292 => X"43",  -- 67
        18293 => X"45",  -- 69
        18294 => X"59",  -- 89
        18295 => X"6A",  -- 106
        18296 => X"82",  -- 130
        18297 => X"8B",  -- 139
        18298 => X"77",  -- 119
        18299 => X"6D",  -- 109
        18300 => X"50",  -- 80
        18301 => X"75",  -- 117
        18302 => X"6A",  -- 106
        18303 => X"68",  -- 104
        18304 => X"88",  -- 136
        18305 => X"77",  -- 119
        18306 => X"46",  -- 70
        18307 => X"20",  -- 32
        18308 => X"2D",  -- 45
        18309 => X"36",  -- 54
        18310 => X"51",  -- 81
        18311 => X"44",  -- 68
        18312 => X"60",  -- 96
        18313 => X"76",  -- 118
        18314 => X"98",  -- 152
        18315 => X"87",  -- 135
        18316 => X"98",  -- 152
        18317 => X"92",  -- 146
        18318 => X"A3",  -- 163
        18319 => X"98",  -- 152
        18320 => X"8F",  -- 143
        18321 => X"94",  -- 148
        18322 => X"95",  -- 149
        18323 => X"8F",  -- 143
        18324 => X"85",  -- 133
        18325 => X"72",  -- 114
        18326 => X"53",  -- 83
        18327 => X"3A",  -- 58
        18328 => X"4A",  -- 74
        18329 => X"61",  -- 97
        18330 => X"44",  -- 68
        18331 => X"38",  -- 56
        18332 => X"2D",  -- 45
        18333 => X"0E",  -- 14
        18334 => X"0D",  -- 13
        18335 => X"0E",  -- 14
        18336 => X"14",  -- 20
        18337 => X"15",  -- 21
        18338 => X"10",  -- 16
        18339 => X"16",  -- 22
        18340 => X"10",  -- 16
        18341 => X"1E",  -- 30
        18342 => X"19",  -- 25
        18343 => X"21",  -- 33
        18344 => X"42",  -- 66
        18345 => X"38",  -- 56
        18346 => X"2F",  -- 47
        18347 => X"39",  -- 57
        18348 => X"47",  -- 71
        18349 => X"47",  -- 71
        18350 => X"4F",  -- 79
        18351 => X"68",  -- 104
        18352 => X"86",  -- 134
        18353 => X"8E",  -- 142
        18354 => X"8E",  -- 142
        18355 => X"8A",  -- 138
        18356 => X"91",  -- 145
        18357 => X"8A",  -- 138
        18358 => X"73",  -- 115
        18359 => X"62",  -- 98
        18360 => X"5D",  -- 93
        18361 => X"49",  -- 73
        18362 => X"28",  -- 40
        18363 => X"12",  -- 18
        18364 => X"0F",  -- 15
        18365 => X"15",  -- 21
        18366 => X"28",  -- 40
        18367 => X"43",  -- 67
        18368 => X"6F",  -- 111
        18369 => X"7E",  -- 126
        18370 => X"74",  -- 116
        18371 => X"68",  -- 104
        18372 => X"4A",  -- 74
        18373 => X"56",  -- 86
        18374 => X"4F",  -- 79
        18375 => X"48",  -- 72
        18376 => X"43",  -- 67
        18377 => X"24",  -- 36
        18378 => X"27",  -- 39
        18379 => X"25",  -- 37
        18380 => X"2C",  -- 44
        18381 => X"38",  -- 56
        18382 => X"45",  -- 69
        18383 => X"25",  -- 37
        18384 => X"37",  -- 55
        18385 => X"3B",  -- 59
        18386 => X"4C",  -- 76
        18387 => X"65",  -- 101
        18388 => X"5F",  -- 95
        18389 => X"5A",  -- 90
        18390 => X"6A",  -- 106
        18391 => X"8A",  -- 138
        18392 => X"8A",  -- 138
        18393 => X"4C",  -- 76
        18394 => X"70",  -- 112
        18395 => X"7C",  -- 124
        18396 => X"87",  -- 135
        18397 => X"87",  -- 135
        18398 => X"95",  -- 149
        18399 => X"49",  -- 73
        18400 => X"4B",  -- 75
        18401 => X"36",  -- 54
        18402 => X"49",  -- 73
        18403 => X"43",  -- 67
        18404 => X"59",  -- 89
        18405 => X"52",  -- 82
        18406 => X"64",  -- 100
        18407 => X"62",  -- 98
        18408 => X"61",  -- 97
        18409 => X"50",  -- 80
        18410 => X"67",  -- 103
        18411 => X"6D",  -- 109
        18412 => X"76",  -- 118
        18413 => X"65",  -- 101
        18414 => X"3A",  -- 58
        18415 => X"A2",  -- 162
        18416 => X"AF",  -- 175
        18417 => X"96",  -- 150
        18418 => X"83",  -- 131
        18419 => X"83",  -- 131
        18420 => X"88",  -- 136
        18421 => X"87",  -- 135
        18422 => X"82",  -- 130
        18423 => X"81",  -- 129
        18424 => X"7F",  -- 127
        18425 => X"7E",  -- 126
        18426 => X"7C",  -- 124
        18427 => X"79",  -- 121
        18428 => X"76",  -- 118
        18429 => X"73",  -- 115
        18430 => X"73",  -- 115
        18431 => X"73",  -- 115
        18432 => X"7E",  -- 126
        18433 => X"78",  -- 120
        18434 => X"73",  -- 115
        18435 => X"75",  -- 117
        18436 => X"82",  -- 130
        18437 => X"90",  -- 144
        18438 => X"92",  -- 146
        18439 => X"8E",  -- 142
        18440 => X"85",  -- 133
        18441 => X"89",  -- 137
        18442 => X"8D",  -- 141
        18443 => X"8C",  -- 140
        18444 => X"89",  -- 137
        18445 => X"8B",  -- 139
        18446 => X"94",  -- 148
        18447 => X"9C",  -- 156
        18448 => X"A1",  -- 161
        18449 => X"A3",  -- 163
        18450 => X"A4",  -- 164
        18451 => X"A3",  -- 163
        18452 => X"A4",  -- 164
        18453 => X"A7",  -- 167
        18454 => X"AC",  -- 172
        18455 => X"AF",  -- 175
        18456 => X"A0",  -- 160
        18457 => X"A4",  -- 164
        18458 => X"9F",  -- 159
        18459 => X"8E",  -- 142
        18460 => X"79",  -- 121
        18461 => X"78",  -- 120
        18462 => X"8C",  -- 140
        18463 => X"A3",  -- 163
        18464 => X"A4",  -- 164
        18465 => X"A2",  -- 162
        18466 => X"A0",  -- 160
        18467 => X"A2",  -- 162
        18468 => X"A2",  -- 162
        18469 => X"A4",  -- 164
        18470 => X"A2",  -- 162
        18471 => X"9F",  -- 159
        18472 => X"9E",  -- 158
        18473 => X"A1",  -- 161
        18474 => X"9E",  -- 158
        18475 => X"95",  -- 149
        18476 => X"8A",  -- 138
        18477 => X"84",  -- 132
        18478 => X"81",  -- 129
        18479 => X"7C",  -- 124
        18480 => X"73",  -- 115
        18481 => X"72",  -- 114
        18482 => X"7A",  -- 122
        18483 => X"81",  -- 129
        18484 => X"7A",  -- 122
        18485 => X"62",  -- 98
        18486 => X"4E",  -- 78
        18487 => X"44",  -- 68
        18488 => X"3A",  -- 58
        18489 => X"4A",  -- 74
        18490 => X"5F",  -- 95
        18491 => X"6D",  -- 109
        18492 => X"75",  -- 117
        18493 => X"7C",  -- 124
        18494 => X"86",  -- 134
        18495 => X"90",  -- 144
        18496 => X"8A",  -- 138
        18497 => X"8D",  -- 141
        18498 => X"92",  -- 146
        18499 => X"99",  -- 153
        18500 => X"9F",  -- 159
        18501 => X"A3",  -- 163
        18502 => X"A5",  -- 165
        18503 => X"A5",  -- 165
        18504 => X"A3",  -- 163
        18505 => X"A2",  -- 162
        18506 => X"9E",  -- 158
        18507 => X"97",  -- 151
        18508 => X"93",  -- 147
        18509 => X"95",  -- 149
        18510 => X"93",  -- 147
        18511 => X"91",  -- 145
        18512 => X"8E",  -- 142
        18513 => X"8F",  -- 143
        18514 => X"8F",  -- 143
        18515 => X"80",  -- 128
        18516 => X"5E",  -- 94
        18517 => X"38",  -- 56
        18518 => X"20",  -- 32
        18519 => X"19",  -- 25
        18520 => X"23",  -- 35
        18521 => X"31",  -- 49
        18522 => X"4B",  -- 75
        18523 => X"6B",  -- 107
        18524 => X"80",  -- 128
        18525 => X"8A",  -- 138
        18526 => X"8F",  -- 143
        18527 => X"92",  -- 146
        18528 => X"96",  -- 150
        18529 => X"97",  -- 151
        18530 => X"92",  -- 146
        18531 => X"92",  -- 146
        18532 => X"93",  -- 147
        18533 => X"82",  -- 130
        18534 => X"6E",  -- 110
        18535 => X"69",  -- 105
        18536 => X"78",  -- 120
        18537 => X"91",  -- 145
        18538 => X"A0",  -- 160
        18539 => X"A4",  -- 164
        18540 => X"A7",  -- 167
        18541 => X"A8",  -- 168
        18542 => X"A4",  -- 164
        18543 => X"A7",  -- 167
        18544 => X"AC",  -- 172
        18545 => X"AB",  -- 171
        18546 => X"A7",  -- 167
        18547 => X"A2",  -- 162
        18548 => X"A9",  -- 169
        18549 => X"B3",  -- 179
        18550 => X"B2",  -- 178
        18551 => X"AA",  -- 170
        18552 => X"BD",  -- 189
        18553 => X"C4",  -- 196
        18554 => X"C5",  -- 197
        18555 => X"C0",  -- 192
        18556 => X"B7",  -- 183
        18557 => X"A9",  -- 169
        18558 => X"A3",  -- 163
        18559 => X"AD",  -- 173
        18560 => X"87",  -- 135
        18561 => X"86",  -- 134
        18562 => X"84",  -- 132
        18563 => X"7F",  -- 127
        18564 => X"7A",  -- 122
        18565 => X"78",  -- 120
        18566 => X"7A",  -- 122
        18567 => X"7E",  -- 126
        18568 => X"82",  -- 130
        18569 => X"86",  -- 134
        18570 => X"8B",  -- 139
        18571 => X"92",  -- 146
        18572 => X"97",  -- 151
        18573 => X"9A",  -- 154
        18574 => X"9B",  -- 155
        18575 => X"9A",  -- 154
        18576 => X"A2",  -- 162
        18577 => X"A0",  -- 160
        18578 => X"3B",  -- 59
        18579 => X"55",  -- 85
        18580 => X"63",  -- 99
        18581 => X"6B",  -- 107
        18582 => X"62",  -- 98
        18583 => X"5D",  -- 93
        18584 => X"4A",  -- 74
        18585 => X"50",  -- 80
        18586 => X"4E",  -- 78
        18587 => X"44",  -- 68
        18588 => X"41",  -- 65
        18589 => X"4F",  -- 79
        18590 => X"60",  -- 96
        18591 => X"6B",  -- 107
        18592 => X"7F",  -- 127
        18593 => X"95",  -- 149
        18594 => X"80",  -- 128
        18595 => X"6A",  -- 106
        18596 => X"7C",  -- 124
        18597 => X"6D",  -- 109
        18598 => X"58",  -- 88
        18599 => X"63",  -- 99
        18600 => X"6B",  -- 107
        18601 => X"75",  -- 117
        18602 => X"82",  -- 130
        18603 => X"87",  -- 135
        18604 => X"83",  -- 131
        18605 => X"7B",  -- 123
        18606 => X"77",  -- 119
        18607 => X"73",  -- 115
        18608 => X"6B",  -- 107
        18609 => X"7D",  -- 125
        18610 => X"6F",  -- 111
        18611 => X"5B",  -- 91
        18612 => X"47",  -- 71
        18613 => X"38",  -- 56
        18614 => X"45",  -- 69
        18615 => X"52",  -- 82
        18616 => X"5E",  -- 94
        18617 => X"6C",  -- 108
        18618 => X"6D",  -- 109
        18619 => X"67",  -- 103
        18620 => X"3C",  -- 60
        18621 => X"7D",  -- 125
        18622 => X"71",  -- 113
        18623 => X"63",  -- 99
        18624 => X"79",  -- 121
        18625 => X"50",  -- 80
        18626 => X"49",  -- 73
        18627 => X"73",  -- 115
        18628 => X"9A",  -- 154
        18629 => X"97",  -- 151
        18630 => X"AA",  -- 170
        18631 => X"B1",  -- 177
        18632 => X"A6",  -- 166
        18633 => X"AB",  -- 171
        18634 => X"B3",  -- 179
        18635 => X"96",  -- 150
        18636 => X"99",  -- 153
        18637 => X"91",  -- 145
        18638 => X"9E",  -- 158
        18639 => X"95",  -- 149
        18640 => X"94",  -- 148
        18641 => X"94",  -- 148
        18642 => X"8C",  -- 140
        18643 => X"73",  -- 115
        18644 => X"52",  -- 82
        18645 => X"34",  -- 52
        18646 => X"23",  -- 35
        18647 => X"1B",  -- 27
        18648 => X"1F",  -- 31
        18649 => X"2E",  -- 46
        18650 => X"23",  -- 35
        18651 => X"16",  -- 22
        18652 => X"1A",  -- 26
        18653 => X"15",  -- 21
        18654 => X"0A",  -- 10
        18655 => X"09",  -- 9
        18656 => X"11",  -- 17
        18657 => X"17",  -- 23
        18658 => X"0E",  -- 14
        18659 => X"12",  -- 18
        18660 => X"17",  -- 23
        18661 => X"3A",  -- 58
        18662 => X"2F",  -- 47
        18663 => X"15",  -- 21
        18664 => X"2A",  -- 42
        18665 => X"1F",  -- 31
        18666 => X"15",  -- 21
        18667 => X"1E",  -- 30
        18668 => X"29",  -- 41
        18669 => X"19",  -- 25
        18670 => X"1B",  -- 27
        18671 => X"3C",  -- 60
        18672 => X"66",  -- 102
        18673 => X"81",  -- 129
        18674 => X"95",  -- 149
        18675 => X"99",  -- 153
        18676 => X"9B",  -- 155
        18677 => X"99",  -- 153
        18678 => X"99",  -- 153
        18679 => X"9E",  -- 158
        18680 => X"97",  -- 151
        18681 => X"8A",  -- 138
        18682 => X"68",  -- 104
        18683 => X"41",  -- 65
        18684 => X"23",  -- 35
        18685 => X"11",  -- 17
        18686 => X"12",  -- 18
        18687 => X"21",  -- 33
        18688 => X"48",  -- 72
        18689 => X"7A",  -- 122
        18690 => X"7D",  -- 125
        18691 => X"6B",  -- 107
        18692 => X"3D",  -- 61
        18693 => X"53",  -- 83
        18694 => X"47",  -- 71
        18695 => X"3C",  -- 60
        18696 => X"39",  -- 57
        18697 => X"31",  -- 49
        18698 => X"21",  -- 33
        18699 => X"20",  -- 32
        18700 => X"4F",  -- 79
        18701 => X"4C",  -- 76
        18702 => X"3C",  -- 60
        18703 => X"3D",  -- 61
        18704 => X"48",  -- 72
        18705 => X"40",  -- 64
        18706 => X"3A",  -- 58
        18707 => X"58",  -- 88
        18708 => X"5A",  -- 90
        18709 => X"6F",  -- 111
        18710 => X"7F",  -- 127
        18711 => X"9E",  -- 158
        18712 => X"7C",  -- 124
        18713 => X"77",  -- 119
        18714 => X"5D",  -- 93
        18715 => X"60",  -- 96
        18716 => X"8F",  -- 143
        18717 => X"8D",  -- 141
        18718 => X"94",  -- 148
        18719 => X"80",  -- 128
        18720 => X"35",  -- 53
        18721 => X"32",  -- 50
        18722 => X"40",  -- 64
        18723 => X"4B",  -- 75
        18724 => X"65",  -- 101
        18725 => X"5C",  -- 92
        18726 => X"6E",  -- 110
        18727 => X"59",  -- 89
        18728 => X"57",  -- 87
        18729 => X"59",  -- 89
        18730 => X"6B",  -- 107
        18731 => X"5D",  -- 93
        18732 => X"6A",  -- 106
        18733 => X"67",  -- 103
        18734 => X"5E",  -- 94
        18735 => X"AB",  -- 171
        18736 => X"A6",  -- 166
        18737 => X"93",  -- 147
        18738 => X"7F",  -- 127
        18739 => X"7B",  -- 123
        18740 => X"7D",  -- 125
        18741 => X"7D",  -- 125
        18742 => X"79",  -- 121
        18743 => X"7A",  -- 122
        18744 => X"7A",  -- 122
        18745 => X"79",  -- 121
        18746 => X"77",  -- 119
        18747 => X"77",  -- 119
        18748 => X"79",  -- 121
        18749 => X"7A",  -- 122
        18750 => X"7E",  -- 126
        18751 => X"80",  -- 128
        18752 => X"84",  -- 132
        18753 => X"89",  -- 137
        18754 => X"88",  -- 136
        18755 => X"82",  -- 130
        18756 => X"7F",  -- 127
        18757 => X"85",  -- 133
        18758 => X"8F",  -- 143
        18759 => X"96",  -- 150
        18760 => X"96",  -- 150
        18761 => X"9D",  -- 157
        18762 => X"A1",  -- 161
        18763 => X"9B",  -- 155
        18764 => X"93",  -- 147
        18765 => X"8F",  -- 143
        18766 => X"95",  -- 149
        18767 => X"9D",  -- 157
        18768 => X"AA",  -- 170
        18769 => X"A5",  -- 165
        18770 => X"A3",  -- 163
        18771 => X"A5",  -- 165
        18772 => X"AC",  -- 172
        18773 => X"B1",  -- 177
        18774 => X"B3",  -- 179
        18775 => X"B3",  -- 179
        18776 => X"A9",  -- 169
        18777 => X"A6",  -- 166
        18778 => X"A3",  -- 163
        18779 => X"98",  -- 152
        18780 => X"82",  -- 130
        18781 => X"74",  -- 116
        18782 => X"7D",  -- 125
        18783 => X"93",  -- 147
        18784 => X"9D",  -- 157
        18785 => X"A2",  -- 162
        18786 => X"A9",  -- 169
        18787 => X"AD",  -- 173
        18788 => X"AD",  -- 173
        18789 => X"AA",  -- 170
        18790 => X"A6",  -- 166
        18791 => X"A4",  -- 164
        18792 => X"A5",  -- 165
        18793 => X"A3",  -- 163
        18794 => X"A1",  -- 161
        18795 => X"9C",  -- 156
        18796 => X"92",  -- 146
        18797 => X"87",  -- 135
        18798 => X"83",  -- 131
        18799 => X"83",  -- 131
        18800 => X"88",  -- 136
        18801 => X"7F",  -- 127
        18802 => X"78",  -- 120
        18803 => X"72",  -- 114
        18804 => X"6F",  -- 111
        18805 => X"66",  -- 102
        18806 => X"55",  -- 85
        18807 => X"48",  -- 72
        18808 => X"3F",  -- 63
        18809 => X"49",  -- 73
        18810 => X"5B",  -- 91
        18811 => X"6E",  -- 110
        18812 => X"7B",  -- 123
        18813 => X"80",  -- 128
        18814 => X"7F",  -- 127
        18815 => X"7B",  -- 123
        18816 => X"8B",  -- 139
        18817 => X"8C",  -- 140
        18818 => X"92",  -- 146
        18819 => X"98",  -- 152
        18820 => X"9D",  -- 157
        18821 => X"A2",  -- 162
        18822 => X"A5",  -- 165
        18823 => X"A6",  -- 166
        18824 => X"A2",  -- 162
        18825 => X"A1",  -- 161
        18826 => X"9E",  -- 158
        18827 => X"9A",  -- 154
        18828 => X"98",  -- 152
        18829 => X"9A",  -- 154
        18830 => X"97",  -- 151
        18831 => X"92",  -- 146
        18832 => X"92",  -- 146
        18833 => X"9B",  -- 155
        18834 => X"94",  -- 148
        18835 => X"74",  -- 116
        18836 => X"4C",  -- 76
        18837 => X"33",  -- 51
        18838 => X"22",  -- 34
        18839 => X"18",  -- 24
        18840 => X"1F",  -- 31
        18841 => X"2E",  -- 46
        18842 => X"4B",  -- 75
        18843 => X"6C",  -- 108
        18844 => X"82",  -- 130
        18845 => X"89",  -- 137
        18846 => X"88",  -- 136
        18847 => X"86",  -- 134
        18848 => X"8C",  -- 140
        18849 => X"8F",  -- 143
        18850 => X"8C",  -- 140
        18851 => X"8C",  -- 140
        18852 => X"8B",  -- 139
        18853 => X"79",  -- 121
        18854 => X"68",  -- 104
        18855 => X"67",  -- 103
        18856 => X"7F",  -- 127
        18857 => X"96",  -- 150
        18858 => X"A2",  -- 162
        18859 => X"A4",  -- 164
        18860 => X"A7",  -- 167
        18861 => X"A6",  -- 166
        18862 => X"A0",  -- 160
        18863 => X"A0",  -- 160
        18864 => X"AD",  -- 173
        18865 => X"AD",  -- 173
        18866 => X"AB",  -- 171
        18867 => X"A9",  -- 169
        18868 => X"AF",  -- 175
        18869 => X"B8",  -- 184
        18870 => X"BB",  -- 187
        18871 => X"B4",  -- 180
        18872 => X"BA",  -- 186
        18873 => X"C4",  -- 196
        18874 => X"C5",  -- 197
        18875 => X"BA",  -- 186
        18876 => X"AC",  -- 172
        18877 => X"9E",  -- 158
        18878 => X"9C",  -- 156
        18879 => X"AA",  -- 170
        18880 => X"88",  -- 136
        18881 => X"87",  -- 135
        18882 => X"86",  -- 134
        18883 => X"82",  -- 130
        18884 => X"7F",  -- 127
        18885 => X"7C",  -- 124
        18886 => X"7E",  -- 126
        18887 => X"80",  -- 128
        18888 => X"84",  -- 132
        18889 => X"88",  -- 136
        18890 => X"8D",  -- 141
        18891 => X"93",  -- 147
        18892 => X"98",  -- 152
        18893 => X"99",  -- 153
        18894 => X"9A",  -- 154
        18895 => X"99",  -- 153
        18896 => X"9D",  -- 157
        18897 => X"9C",  -- 156
        18898 => X"56",  -- 86
        18899 => X"3D",  -- 61
        18900 => X"5E",  -- 94
        18901 => X"60",  -- 96
        18902 => X"5E",  -- 94
        18903 => X"42",  -- 66
        18904 => X"3F",  -- 63
        18905 => X"48",  -- 72
        18906 => X"4D",  -- 77
        18907 => X"4B",  -- 75
        18908 => X"4A",  -- 74
        18909 => X"53",  -- 83
        18910 => X"5E",  -- 94
        18911 => X"67",  -- 103
        18912 => X"82",  -- 130
        18913 => X"80",  -- 128
        18914 => X"68",  -- 104
        18915 => X"58",  -- 88
        18916 => X"84",  -- 132
        18917 => X"75",  -- 117
        18918 => X"73",  -- 115
        18919 => X"8F",  -- 143
        18920 => X"90",  -- 144
        18921 => X"85",  -- 133
        18922 => X"70",  -- 112
        18923 => X"63",  -- 99
        18924 => X"6A",  -- 106
        18925 => X"7B",  -- 123
        18926 => X"89",  -- 137
        18927 => X"93",  -- 147
        18928 => X"70",  -- 112
        18929 => X"70",  -- 112
        18930 => X"65",  -- 101
        18931 => X"65",  -- 101
        18932 => X"57",  -- 87
        18933 => X"3F",  -- 63
        18934 => X"43",  -- 67
        18935 => X"4E",  -- 78
        18936 => X"4C",  -- 76
        18937 => X"4E",  -- 78
        18938 => X"52",  -- 82
        18939 => X"47",  -- 71
        18940 => X"32",  -- 50
        18941 => X"6A",  -- 106
        18942 => X"67",  -- 103
        18943 => X"6C",  -- 108
        18944 => X"68",  -- 104
        18945 => X"50",  -- 80
        18946 => X"6E",  -- 110
        18947 => X"AE",  -- 174
        18948 => X"C3",  -- 195
        18949 => X"B3",  -- 179
        18950 => X"C1",  -- 193
        18951 => X"D1",  -- 209
        18952 => X"C3",  -- 195
        18953 => X"B8",  -- 184
        18954 => X"B2",  -- 178
        18955 => X"9E",  -- 158
        18956 => X"A9",  -- 169
        18957 => X"A1",  -- 161
        18958 => X"9D",  -- 157
        18959 => X"88",  -- 136
        18960 => X"83",  -- 131
        18961 => X"72",  -- 114
        18962 => X"58",  -- 88
        18963 => X"38",  -- 56
        18964 => X"19",  -- 25
        18965 => X"09",  -- 9
        18966 => X"0E",  -- 14
        18967 => X"18",  -- 24
        18968 => X"0A",  -- 10
        18969 => X"12",  -- 18
        18970 => X"1D",  -- 29
        18971 => X"1C",  -- 28
        18972 => X"34",  -- 52
        18973 => X"3F",  -- 63
        18974 => X"19",  -- 25
        18975 => X"08",  -- 8
        18976 => X"0C",  -- 12
        18977 => X"14",  -- 20
        18978 => X"0D",  -- 13
        18979 => X"1F",  -- 31
        18980 => X"33",  -- 51
        18981 => X"5F",  -- 95
        18982 => X"66",  -- 102
        18983 => X"4C",  -- 76
        18984 => X"27",  -- 39
        18985 => X"15",  -- 21
        18986 => X"0F",  -- 15
        18987 => X"17",  -- 23
        18988 => X"19",  -- 25
        18989 => X"11",  -- 17
        18990 => X"0D",  -- 13
        18991 => X"13",  -- 19
        18992 => X"32",  -- 50
        18993 => X"57",  -- 87
        18994 => X"79",  -- 121
        18995 => X"8A",  -- 138
        18996 => X"92",  -- 146
        18997 => X"93",  -- 147
        18998 => X"9A",  -- 154
        18999 => X"A9",  -- 169
        19000 => X"B6",  -- 182
        19001 => X"AE",  -- 174
        19002 => X"A0",  -- 160
        19003 => X"8F",  -- 143
        19004 => X"6D",  -- 109
        19005 => X"3A",  -- 58
        19006 => X"1B",  -- 27
        19007 => X"1D",  -- 29
        19008 => X"1C",  -- 28
        19009 => X"51",  -- 81
        19010 => X"64",  -- 100
        19011 => X"56",  -- 86
        19012 => X"37",  -- 55
        19013 => X"3C",  -- 60
        19014 => X"30",  -- 48
        19015 => X"2B",  -- 43
        19016 => X"35",  -- 53
        19017 => X"1E",  -- 30
        19018 => X"25",  -- 37
        19019 => X"33",  -- 51
        19020 => X"46",  -- 70
        19021 => X"3A",  -- 58
        19022 => X"3F",  -- 63
        19023 => X"3E",  -- 62
        19024 => X"57",  -- 87
        19025 => X"47",  -- 71
        19026 => X"32",  -- 50
        19027 => X"4D",  -- 77
        19028 => X"3E",  -- 62
        19029 => X"50",  -- 80
        19030 => X"5E",  -- 94
        19031 => X"89",  -- 137
        19032 => X"8F",  -- 143
        19033 => X"83",  -- 131
        19034 => X"64",  -- 100
        19035 => X"69",  -- 105
        19036 => X"65",  -- 101
        19037 => X"83",  -- 131
        19038 => X"AE",  -- 174
        19039 => X"73",  -- 115
        19040 => X"27",  -- 39
        19041 => X"26",  -- 38
        19042 => X"38",  -- 56
        19043 => X"42",  -- 66
        19044 => X"5B",  -- 91
        19045 => X"5F",  -- 95
        19046 => X"65",  -- 101
        19047 => X"4D",  -- 77
        19048 => X"4E",  -- 78
        19049 => X"60",  -- 96
        19050 => X"67",  -- 103
        19051 => X"5F",  -- 95
        19052 => X"67",  -- 103
        19053 => X"53",  -- 83
        19054 => X"9C",  -- 156
        19055 => X"BC",  -- 188
        19056 => X"B1",  -- 177
        19057 => X"9B",  -- 155
        19058 => X"85",  -- 133
        19059 => X"79",  -- 121
        19060 => X"77",  -- 119
        19061 => X"79",  -- 121
        19062 => X"7A",  -- 122
        19063 => X"7F",  -- 127
        19064 => X"76",  -- 118
        19065 => X"75",  -- 117
        19066 => X"76",  -- 118
        19067 => X"79",  -- 121
        19068 => X"7B",  -- 123
        19069 => X"80",  -- 128
        19070 => X"84",  -- 132
        19071 => X"85",  -- 133
        19072 => X"82",  -- 130
        19073 => X"89",  -- 137
        19074 => X"8E",  -- 142
        19075 => X"8A",  -- 138
        19076 => X"82",  -- 130
        19077 => X"81",  -- 129
        19078 => X"89",  -- 137
        19079 => X"90",  -- 144
        19080 => X"A3",  -- 163
        19081 => X"A4",  -- 164
        19082 => X"A4",  -- 164
        19083 => X"A6",  -- 166
        19084 => X"A7",  -- 167
        19085 => X"A5",  -- 165
        19086 => X"A3",  -- 163
        19087 => X"A2",  -- 162
        19088 => X"AC",  -- 172
        19089 => X"AB",  -- 171
        19090 => X"AE",  -- 174
        19091 => X"B3",  -- 179
        19092 => X"B9",  -- 185
        19093 => X"BA",  -- 186
        19094 => X"B6",  -- 182
        19095 => X"B1",  -- 177
        19096 => X"B1",  -- 177
        19097 => X"AC",  -- 172
        19098 => X"A6",  -- 166
        19099 => X"9A",  -- 154
        19100 => X"83",  -- 131
        19101 => X"71",  -- 113
        19102 => X"76",  -- 118
        19103 => X"87",  -- 135
        19104 => X"9B",  -- 155
        19105 => X"A5",  -- 165
        19106 => X"AE",  -- 174
        19107 => X"B2",  -- 178
        19108 => X"B0",  -- 176
        19109 => X"AC",  -- 172
        19110 => X"A8",  -- 168
        19111 => X"A6",  -- 166
        19112 => X"AA",  -- 170
        19113 => X"A6",  -- 166
        19114 => X"A3",  -- 163
        19115 => X"A0",  -- 160
        19116 => X"95",  -- 149
        19117 => X"88",  -- 136
        19118 => X"86",  -- 134
        19119 => X"8C",  -- 140
        19120 => X"8B",  -- 139
        19121 => X"89",  -- 137
        19122 => X"83",  -- 131
        19123 => X"80",  -- 128
        19124 => X"7F",  -- 127
        19125 => X"74",  -- 116
        19126 => X"59",  -- 89
        19127 => X"3D",  -- 61
        19128 => X"37",  -- 55
        19129 => X"43",  -- 67
        19130 => X"56",  -- 86
        19131 => X"6E",  -- 110
        19132 => X"82",  -- 130
        19133 => X"88",  -- 136
        19134 => X"86",  -- 134
        19135 => X"80",  -- 128
        19136 => X"89",  -- 137
        19137 => X"8B",  -- 139
        19138 => X"91",  -- 145
        19139 => X"96",  -- 150
        19140 => X"9C",  -- 156
        19141 => X"A1",  -- 161
        19142 => X"A8",  -- 168
        19143 => X"AB",  -- 171
        19144 => X"A8",  -- 168
        19145 => X"A7",  -- 167
        19146 => X"A4",  -- 164
        19147 => X"A1",  -- 161
        19148 => X"A1",  -- 161
        19149 => X"A2",  -- 162
        19150 => X"9D",  -- 157
        19151 => X"95",  -- 149
        19152 => X"9C",  -- 156
        19153 => X"9E",  -- 158
        19154 => X"8E",  -- 142
        19155 => X"6A",  -- 106
        19156 => X"47",  -- 71
        19157 => X"30",  -- 48
        19158 => X"24",  -- 36
        19159 => X"1A",  -- 26
        19160 => X"1B",  -- 27
        19161 => X"30",  -- 48
        19162 => X"50",  -- 80
        19163 => X"6F",  -- 111
        19164 => X"81",  -- 129
        19165 => X"87",  -- 135
        19166 => X"84",  -- 132
        19167 => X"82",  -- 130
        19168 => X"84",  -- 132
        19169 => X"89",  -- 137
        19170 => X"8B",  -- 139
        19171 => X"8E",  -- 142
        19172 => X"89",  -- 137
        19173 => X"78",  -- 120
        19174 => X"68",  -- 104
        19175 => X"6A",  -- 106
        19176 => X"85",  -- 133
        19177 => X"9B",  -- 155
        19178 => X"A8",  -- 168
        19179 => X"AA",  -- 170
        19180 => X"AE",  -- 174
        19181 => X"AC",  -- 172
        19182 => X"A6",  -- 166
        19183 => X"A5",  -- 165
        19184 => X"A3",  -- 163
        19185 => X"A5",  -- 165
        19186 => X"A5",  -- 165
        19187 => X"A4",  -- 164
        19188 => X"A9",  -- 169
        19189 => X"B2",  -- 178
        19190 => X"B2",  -- 178
        19191 => X"AF",  -- 175
        19192 => X"B4",  -- 180
        19193 => X"C0",  -- 192
        19194 => X"C1",  -- 193
        19195 => X"B7",  -- 183
        19196 => X"AB",  -- 171
        19197 => X"9F",  -- 159
        19198 => X"9E",  -- 158
        19199 => X"AA",  -- 170
        19200 => X"92",  -- 146
        19201 => X"91",  -- 145
        19202 => X"8E",  -- 142
        19203 => X"8C",  -- 140
        19204 => X"8A",  -- 138
        19205 => X"89",  -- 137
        19206 => X"8A",  -- 138
        19207 => X"8C",  -- 140
        19208 => X"90",  -- 144
        19209 => X"92",  -- 146
        19210 => X"94",  -- 148
        19211 => X"97",  -- 151
        19212 => X"9A",  -- 154
        19213 => X"9B",  -- 155
        19214 => X"9B",  -- 155
        19215 => X"9B",  -- 155
        19216 => X"A9",  -- 169
        19217 => X"97",  -- 151
        19218 => X"78",  -- 120
        19219 => X"3C",  -- 60
        19220 => X"52",  -- 82
        19221 => X"51",  -- 81
        19222 => X"56",  -- 86
        19223 => X"4E",  -- 78
        19224 => X"42",  -- 66
        19225 => X"47",  -- 71
        19226 => X"4B",  -- 75
        19227 => X"4B",  -- 75
        19228 => X"4C",  -- 76
        19229 => X"52",  -- 82
        19230 => X"58",  -- 88
        19231 => X"5C",  -- 92
        19232 => X"61",  -- 97
        19233 => X"4A",  -- 74
        19234 => X"4D",  -- 77
        19235 => X"85",  -- 133
        19236 => X"65",  -- 101
        19237 => X"8B",  -- 139
        19238 => X"84",  -- 132
        19239 => X"73",  -- 115
        19240 => X"5C",  -- 92
        19241 => X"59",  -- 89
        19242 => X"48",  -- 72
        19243 => X"42",  -- 66
        19244 => X"54",  -- 84
        19245 => X"65",  -- 101
        19246 => X"71",  -- 113
        19247 => X"7D",  -- 125
        19248 => X"88",  -- 136
        19249 => X"75",  -- 117
        19250 => X"63",  -- 99
        19251 => X"6B",  -- 107
        19252 => X"5D",  -- 93
        19253 => X"43",  -- 67
        19254 => X"4D",  -- 77
        19255 => X"5E",  -- 94
        19256 => X"56",  -- 86
        19257 => X"4A",  -- 74
        19258 => X"42",  -- 66
        19259 => X"2F",  -- 47
        19260 => X"31",  -- 49
        19261 => X"3B",  -- 59
        19262 => X"4A",  -- 74
        19263 => X"76",  -- 118
        19264 => X"72",  -- 114
        19265 => X"8A",  -- 138
        19266 => X"B6",  -- 182
        19267 => X"CC",  -- 204
        19268 => X"C2",  -- 194
        19269 => X"C8",  -- 200
        19270 => X"C6",  -- 198
        19271 => X"BC",  -- 188
        19272 => X"C0",  -- 192
        19273 => X"B4",  -- 180
        19274 => X"AA",  -- 170
        19275 => X"9F",  -- 159
        19276 => X"A9",  -- 169
        19277 => X"A3",  -- 163
        19278 => X"99",  -- 153
        19279 => X"82",  -- 130
        19280 => X"51",  -- 81
        19281 => X"39",  -- 57
        19282 => X"1E",  -- 30
        19283 => X"14",  -- 20
        19284 => X"15",  -- 21
        19285 => X"14",  -- 20
        19286 => X"10",  -- 16
        19287 => X"0C",  -- 12
        19288 => X"0F",  -- 15
        19289 => X"0A",  -- 10
        19290 => X"1D",  -- 29
        19291 => X"26",  -- 38
        19292 => X"49",  -- 73
        19293 => X"5E",  -- 94
        19294 => X"29",  -- 41
        19295 => X"09",  -- 9
        19296 => X"0C",  -- 12
        19297 => X"18",  -- 24
        19298 => X"1D",  -- 29
        19299 => X"49",  -- 73
        19300 => X"61",  -- 97
        19301 => X"7F",  -- 127
        19302 => X"90",  -- 144
        19303 => X"8B",  -- 139
        19304 => X"46",  -- 70
        19305 => X"16",  -- 22
        19306 => X"09",  -- 9
        19307 => X"11",  -- 17
        19308 => X"0F",  -- 15
        19309 => X"15",  -- 21
        19310 => X"19",  -- 25
        19311 => X"05",  -- 5
        19312 => X"12",  -- 18
        19313 => X"25",  -- 37
        19314 => X"41",  -- 65
        19315 => X"64",  -- 100
        19316 => X"87",  -- 135
        19317 => X"95",  -- 149
        19318 => X"96",  -- 150
        19319 => X"9A",  -- 154
        19320 => X"BB",  -- 187
        19321 => X"B5",  -- 181
        19322 => X"B2",  -- 178
        19323 => X"B9",  -- 185
        19324 => X"B4",  -- 180
        19325 => X"88",  -- 136
        19326 => X"56",  -- 86
        19327 => X"3D",  -- 61
        19328 => X"2A",  -- 42
        19329 => X"42",  -- 66
        19330 => X"56",  -- 86
        19331 => X"47",  -- 71
        19332 => X"42",  -- 66
        19333 => X"26",  -- 38
        19334 => X"26",  -- 38
        19335 => X"2B",  -- 43
        19336 => X"23",  -- 35
        19337 => X"39",  -- 57
        19338 => X"2F",  -- 47
        19339 => X"29",  -- 41
        19340 => X"59",  -- 89
        19341 => X"43",  -- 67
        19342 => X"33",  -- 51
        19343 => X"51",  -- 81
        19344 => X"4B",  -- 75
        19345 => X"41",  -- 65
        19346 => X"35",  -- 53
        19347 => X"4E",  -- 78
        19348 => X"2A",  -- 42
        19349 => X"24",  -- 36
        19350 => X"2D",  -- 45
        19351 => X"60",  -- 96
        19352 => X"7A",  -- 122
        19353 => X"87",  -- 135
        19354 => X"79",  -- 121
        19355 => X"71",  -- 113
        19356 => X"3C",  -- 60
        19357 => X"64",  -- 100
        19358 => X"AB",  -- 171
        19359 => X"62",  -- 98
        19360 => X"21",  -- 33
        19361 => X"1C",  -- 28
        19362 => X"3E",  -- 62
        19363 => X"34",  -- 52
        19364 => X"3D",  -- 61
        19365 => X"4F",  -- 79
        19366 => X"4B",  -- 75
        19367 => X"4B",  -- 75
        19368 => X"53",  -- 83
        19369 => X"5D",  -- 93
        19370 => X"63",  -- 99
        19371 => X"71",  -- 113
        19372 => X"57",  -- 87
        19373 => X"58",  -- 88
        19374 => X"B2",  -- 178
        19375 => X"C8",  -- 200
        19376 => X"B7",  -- 183
        19377 => X"A2",  -- 162
        19378 => X"8B",  -- 139
        19379 => X"7C",  -- 124
        19380 => X"78",  -- 120
        19381 => X"77",  -- 119
        19382 => X"79",  -- 121
        19383 => X"7D",  -- 125
        19384 => X"7A",  -- 122
        19385 => X"79",  -- 121
        19386 => X"79",  -- 121
        19387 => X"7C",  -- 124
        19388 => X"7D",  -- 125
        19389 => X"7E",  -- 126
        19390 => X"7F",  -- 127
        19391 => X"7C",  -- 124
        19392 => X"85",  -- 133
        19393 => X"81",  -- 129
        19394 => X"81",  -- 129
        19395 => X"88",  -- 136
        19396 => X"91",  -- 145
        19397 => X"93",  -- 147
        19398 => X"8B",  -- 139
        19399 => X"85",  -- 133
        19400 => X"93",  -- 147
        19401 => X"94",  -- 148
        19402 => X"9A",  -- 154
        19403 => X"A2",  -- 162
        19404 => X"A9",  -- 169
        19405 => X"AB",  -- 171
        19406 => X"A8",  -- 168
        19407 => X"A3",  -- 163
        19408 => X"A8",  -- 168
        19409 => X"AE",  -- 174
        19410 => X"B6",  -- 182
        19411 => X"BD",  -- 189
        19412 => X"BF",  -- 191
        19413 => X"BD",  -- 189
        19414 => X"B8",  -- 184
        19415 => X"B5",  -- 181
        19416 => X"AD",  -- 173
        19417 => X"AF",  -- 175
        19418 => X"A8",  -- 168
        19419 => X"97",  -- 151
        19420 => X"84",  -- 132
        19421 => X"7D",  -- 125
        19422 => X"84",  -- 132
        19423 => X"8C",  -- 140
        19424 => X"A1",  -- 161
        19425 => X"A9",  -- 169
        19426 => X"B2",  -- 178
        19427 => X"B6",  -- 182
        19428 => X"B2",  -- 178
        19429 => X"AC",  -- 172
        19430 => X"A9",  -- 169
        19431 => X"AA",  -- 170
        19432 => X"B0",  -- 176
        19433 => X"AA",  -- 170
        19434 => X"A5",  -- 165
        19435 => X"A1",  -- 161
        19436 => X"98",  -- 152
        19437 => X"8C",  -- 140
        19438 => X"8D",  -- 141
        19439 => X"94",  -- 148
        19440 => X"92",  -- 146
        19441 => X"90",  -- 144
        19442 => X"89",  -- 137
        19443 => X"84",  -- 132
        19444 => X"82",  -- 130
        19445 => X"76",  -- 118
        19446 => X"54",  -- 84
        19447 => X"34",  -- 52
        19448 => X"28",  -- 40
        19449 => X"40",  -- 64
        19450 => X"60",  -- 96
        19451 => X"72",  -- 114
        19452 => X"77",  -- 119
        19453 => X"7B",  -- 123
        19454 => X"86",  -- 134
        19455 => X"90",  -- 144
        19456 => X"89",  -- 137
        19457 => X"8C",  -- 140
        19458 => X"8F",  -- 143
        19459 => X"93",  -- 147
        19460 => X"99",  -- 153
        19461 => X"9D",  -- 157
        19462 => X"A4",  -- 164
        19463 => X"A9",  -- 169
        19464 => X"AC",  -- 172
        19465 => X"AB",  -- 171
        19466 => X"A7",  -- 167
        19467 => X"A6",  -- 166
        19468 => X"A6",  -- 166
        19469 => X"A9",  -- 169
        19470 => X"A4",  -- 164
        19471 => X"9B",  -- 155
        19472 => X"9D",  -- 157
        19473 => X"94",  -- 148
        19474 => X"81",  -- 129
        19475 => X"69",  -- 105
        19476 => X"4E",  -- 78
        19477 => X"33",  -- 51
        19478 => X"1F",  -- 31
        19479 => X"17",  -- 23
        19480 => X"1F",  -- 31
        19481 => X"3A",  -- 58
        19482 => X"5E",  -- 94
        19483 => X"79",  -- 121
        19484 => X"84",  -- 132
        19485 => X"87",  -- 135
        19486 => X"87",  -- 135
        19487 => X"88",  -- 136
        19488 => X"8A",  -- 138
        19489 => X"90",  -- 144
        19490 => X"94",  -- 148
        19491 => X"95",  -- 149
        19492 => X"8E",  -- 142
        19493 => X"7A",  -- 122
        19494 => X"6D",  -- 109
        19495 => X"74",  -- 116
        19496 => X"87",  -- 135
        19497 => X"9C",  -- 156
        19498 => X"A8",  -- 168
        19499 => X"AA",  -- 170
        19500 => X"B2",  -- 178
        19501 => X"B2",  -- 178
        19502 => X"AA",  -- 170
        19503 => X"A7",  -- 167
        19504 => X"9E",  -- 158
        19505 => X"9E",  -- 158
        19506 => X"A0",  -- 160
        19507 => X"A3",  -- 163
        19508 => X"A7",  -- 167
        19509 => X"AC",  -- 172
        19510 => X"AC",  -- 172
        19511 => X"A9",  -- 169
        19512 => X"B2",  -- 178
        19513 => X"BF",  -- 191
        19514 => X"C2",  -- 194
        19515 => X"BC",  -- 188
        19516 => X"B6",  -- 182
        19517 => X"AB",  -- 171
        19518 => X"A6",  -- 166
        19519 => X"AB",  -- 171
        19520 => X"A0",  -- 160
        19521 => X"9E",  -- 158
        19522 => X"9D",  -- 157
        19523 => X"9A",  -- 154
        19524 => X"9A",  -- 154
        19525 => X"9A",  -- 154
        19526 => X"9A",  -- 154
        19527 => X"9B",  -- 155
        19528 => X"9A",  -- 154
        19529 => X"9B",  -- 155
        19530 => X"9B",  -- 155
        19531 => X"9A",  -- 154
        19532 => X"9C",  -- 156
        19533 => X"9B",  -- 155
        19534 => X"9C",  -- 156
        19535 => X"9B",  -- 155
        19536 => X"9D",  -- 157
        19537 => X"98",  -- 152
        19538 => X"8A",  -- 138
        19539 => X"47",  -- 71
        19540 => X"2C",  -- 44
        19541 => X"4A",  -- 74
        19542 => X"4F",  -- 79
        19543 => X"51",  -- 81
        19544 => X"4B",  -- 75
        19545 => X"49",  -- 73
        19546 => X"44",  -- 68
        19547 => X"40",  -- 64
        19548 => X"41",  -- 65
        19549 => X"44",  -- 68
        19550 => X"4A",  -- 74
        19551 => X"4E",  -- 78
        19552 => X"3E",  -- 62
        19553 => X"2A",  -- 42
        19554 => X"61",  -- 97
        19555 => X"52",  -- 82
        19556 => X"68",  -- 104
        19557 => X"54",  -- 84
        19558 => X"68",  -- 104
        19559 => X"2A",  -- 42
        19560 => X"2A",  -- 42
        19561 => X"3A",  -- 58
        19562 => X"3B",  -- 59
        19563 => X"3B",  -- 59
        19564 => X"46",  -- 70
        19565 => X"44",  -- 68
        19566 => X"41",  -- 65
        19567 => X"4F",  -- 79
        19568 => X"61",  -- 97
        19569 => X"58",  -- 88
        19570 => X"56",  -- 86
        19571 => X"66",  -- 102
        19572 => X"57",  -- 87
        19573 => X"43",  -- 67
        19574 => X"55",  -- 85
        19575 => X"65",  -- 101
        19576 => X"51",  -- 81
        19577 => X"46",  -- 70
        19578 => X"3A",  -- 58
        19579 => X"33",  -- 51
        19580 => X"44",  -- 68
        19581 => X"2D",  -- 45
        19582 => X"4D",  -- 77
        19583 => X"8A",  -- 138
        19584 => X"8F",  -- 143
        19585 => X"A3",  -- 163
        19586 => X"B9",  -- 185
        19587 => X"B5",  -- 181
        19588 => X"9D",  -- 157
        19589 => X"A0",  -- 160
        19590 => X"90",  -- 144
        19591 => X"89",  -- 137
        19592 => X"A2",  -- 162
        19593 => X"A4",  -- 164
        19594 => X"A6",  -- 166
        19595 => X"9C",  -- 156
        19596 => X"90",  -- 144
        19597 => X"75",  -- 117
        19598 => X"5D",  -- 93
        19599 => X"4B",  -- 75
        19600 => X"20",  -- 32
        19601 => X"18",  -- 24
        19602 => X"13",  -- 19
        19603 => X"15",  -- 21
        19604 => X"1D",  -- 29
        19605 => X"20",  -- 32
        19606 => X"17",  -- 23
        19607 => X"0E",  -- 14
        19608 => X"17",  -- 23
        19609 => X"08",  -- 8
        19610 => X"13",  -- 19
        19611 => X"20",  -- 32
        19612 => X"48",  -- 72
        19613 => X"65",  -- 101
        19614 => X"41",  -- 65
        19615 => X"20",  -- 32
        19616 => X"1D",  -- 29
        19617 => X"3A",  -- 58
        19618 => X"43",  -- 67
        19619 => X"76",  -- 118
        19620 => X"88",  -- 136
        19621 => X"86",  -- 134
        19622 => X"8C",  -- 140
        19623 => X"95",  -- 149
        19624 => X"7E",  -- 126
        19625 => X"36",  -- 54
        19626 => X"15",  -- 21
        19627 => X"15",  -- 21
        19628 => X"09",  -- 9
        19629 => X"0C",  -- 12
        19630 => X"16",  -- 22
        19631 => X"0C",  -- 12
        19632 => X"08",  -- 8
        19633 => X"0E",  -- 14
        19634 => X"17",  -- 23
        19635 => X"2F",  -- 47
        19636 => X"53",  -- 83
        19637 => X"71",  -- 113
        19638 => X"8A",  -- 138
        19639 => X"A4",  -- 164
        19640 => X"A4",  -- 164
        19641 => X"B7",  -- 183
        19642 => X"BB",  -- 187
        19643 => X"B9",  -- 185
        19644 => X"BF",  -- 191
        19645 => X"B9",  -- 185
        19646 => X"9A",  -- 154
        19647 => X"80",  -- 128
        19648 => X"77",  -- 119
        19649 => X"6A",  -- 106
        19650 => X"65",  -- 101
        19651 => X"48",  -- 72
        19652 => X"4E",  -- 78
        19653 => X"1F",  -- 31
        19654 => X"1F",  -- 31
        19655 => X"2A",  -- 42
        19656 => X"2A",  -- 42
        19657 => X"35",  -- 53
        19658 => X"44",  -- 68
        19659 => X"3E",  -- 62
        19660 => X"54",  -- 84
        19661 => X"5F",  -- 95
        19662 => X"66",  -- 102
        19663 => X"56",  -- 86
        19664 => X"4E",  -- 78
        19665 => X"33",  -- 51
        19666 => X"21",  -- 33
        19667 => X"3C",  -- 60
        19668 => X"2E",  -- 46
        19669 => X"29",  -- 41
        19670 => X"28",  -- 40
        19671 => X"47",  -- 71
        19672 => X"4F",  -- 79
        19673 => X"81",  -- 129
        19674 => X"84",  -- 132
        19675 => X"6E",  -- 110
        19676 => X"3E",  -- 62
        19677 => X"4C",  -- 76
        19678 => X"8C",  -- 140
        19679 => X"69",  -- 105
        19680 => X"28",  -- 40
        19681 => X"25",  -- 37
        19682 => X"4C",  -- 76
        19683 => X"34",  -- 52
        19684 => X"2A",  -- 42
        19685 => X"3D",  -- 61
        19686 => X"3D",  -- 61
        19687 => X"53",  -- 83
        19688 => X"5B",  -- 91
        19689 => X"64",  -- 100
        19690 => X"61",  -- 97
        19691 => X"55",  -- 85
        19692 => X"34",  -- 52
        19693 => X"90",  -- 144
        19694 => X"B8",  -- 184
        19695 => X"C7",  -- 199
        19696 => X"B0",  -- 176
        19697 => X"9F",  -- 159
        19698 => X"8B",  -- 139
        19699 => X"7D",  -- 125
        19700 => X"79",  -- 121
        19701 => X"76",  -- 118
        19702 => X"72",  -- 114
        19703 => X"6F",  -- 111
        19704 => X"7B",  -- 123
        19705 => X"7A",  -- 122
        19706 => X"7B",  -- 123
        19707 => X"7F",  -- 127
        19708 => X"83",  -- 131
        19709 => X"86",  -- 134
        19710 => X"83",  -- 131
        19711 => X"82",  -- 130
        19712 => X"85",  -- 133
        19713 => X"85",  -- 133
        19714 => X"89",  -- 137
        19715 => X"8F",  -- 143
        19716 => X"90",  -- 144
        19717 => X"8C",  -- 140
        19718 => X"88",  -- 136
        19719 => X"83",  -- 131
        19720 => X"89",  -- 137
        19721 => X"92",  -- 146
        19722 => X"9D",  -- 157
        19723 => X"A3",  -- 163
        19724 => X"A4",  -- 164
        19725 => X"A5",  -- 165
        19726 => X"A8",  -- 168
        19727 => X"AC",  -- 172
        19728 => X"B0",  -- 176
        19729 => X"B5",  -- 181
        19730 => X"BB",  -- 187
        19731 => X"BB",  -- 187
        19732 => X"B8",  -- 184
        19733 => X"B5",  -- 181
        19734 => X"B4",  -- 180
        19735 => X"B5",  -- 181
        19736 => X"AD",  -- 173
        19737 => X"B2",  -- 178
        19738 => X"AB",  -- 171
        19739 => X"98",  -- 152
        19740 => X"83",  -- 131
        19741 => X"7D",  -- 125
        19742 => X"85",  -- 133
        19743 => X"8D",  -- 141
        19744 => X"A7",  -- 167
        19745 => X"AD",  -- 173
        19746 => X"B4",  -- 180
        19747 => X"B5",  -- 181
        19748 => X"B2",  -- 178
        19749 => X"AF",  -- 175
        19750 => X"AC",  -- 172
        19751 => X"AD",  -- 173
        19752 => X"AE",  -- 174
        19753 => X"A9",  -- 169
        19754 => X"A4",  -- 164
        19755 => X"9E",  -- 158
        19756 => X"98",  -- 152
        19757 => X"92",  -- 146
        19758 => X"92",  -- 146
        19759 => X"94",  -- 148
        19760 => X"99",  -- 153
        19761 => X"92",  -- 146
        19762 => X"86",  -- 134
        19763 => X"7C",  -- 124
        19764 => X"76",  -- 118
        19765 => X"6A",  -- 106
        19766 => X"50",  -- 80
        19767 => X"35",  -- 53
        19768 => X"2B",  -- 43
        19769 => X"3E",  -- 62
        19770 => X"5C",  -- 92
        19771 => X"70",  -- 112
        19772 => X"7B",  -- 123
        19773 => X"82",  -- 130
        19774 => X"8D",  -- 141
        19775 => X"94",  -- 148
        19776 => X"8D",  -- 141
        19777 => X"90",  -- 144
        19778 => X"91",  -- 145
        19779 => X"93",  -- 147
        19780 => X"94",  -- 148
        19781 => X"96",  -- 150
        19782 => X"9D",  -- 157
        19783 => X"A2",  -- 162
        19784 => X"A8",  -- 168
        19785 => X"A9",  -- 169
        19786 => X"A6",  -- 166
        19787 => X"A4",  -- 164
        19788 => X"A5",  -- 165
        19789 => X"AA",  -- 170
        19790 => X"A7",  -- 167
        19791 => X"A2",  -- 162
        19792 => X"9C",  -- 156
        19793 => X"90",  -- 144
        19794 => X"83",  -- 131
        19795 => X"76",  -- 118
        19796 => X"5A",  -- 90
        19797 => X"35",  -- 53
        19798 => X"1D",  -- 29
        19799 => X"15",  -- 21
        19800 => X"24",  -- 36
        19801 => X"43",  -- 67
        19802 => X"66",  -- 102
        19803 => X"7D",  -- 125
        19804 => X"83",  -- 131
        19805 => X"86",  -- 134
        19806 => X"89",  -- 137
        19807 => X"8C",  -- 140
        19808 => X"89",  -- 137
        19809 => X"8F",  -- 143
        19810 => X"91",  -- 145
        19811 => X"90",  -- 144
        19812 => X"85",  -- 133
        19813 => X"70",  -- 112
        19814 => X"69",  -- 105
        19815 => X"76",  -- 118
        19816 => X"8A",  -- 138
        19817 => X"9B",  -- 155
        19818 => X"A5",  -- 165
        19819 => X"A8",  -- 168
        19820 => X"AE",  -- 174
        19821 => X"AE",  -- 174
        19822 => X"A4",  -- 164
        19823 => X"A1",  -- 161
        19824 => X"98",  -- 152
        19825 => X"9B",  -- 155
        19826 => X"A0",  -- 160
        19827 => X"A9",  -- 169
        19828 => X"B3",  -- 179
        19829 => X"B9",  -- 185
        19830 => X"B7",  -- 183
        19831 => X"B4",  -- 180
        19832 => X"B0",  -- 176
        19833 => X"BD",  -- 189
        19834 => X"C1",  -- 193
        19835 => X"BF",  -- 191
        19836 => X"BC",  -- 188
        19837 => X"B3",  -- 179
        19838 => X"A8",  -- 168
        19839 => X"A6",  -- 166
        19840 => X"A8",  -- 168
        19841 => X"A6",  -- 166
        19842 => X"A5",  -- 165
        19843 => X"A5",  -- 165
        19844 => X"A6",  -- 166
        19845 => X"A6",  -- 166
        19846 => X"A6",  -- 166
        19847 => X"A4",  -- 164
        19848 => X"A0",  -- 160
        19849 => X"A0",  -- 160
        19850 => X"9E",  -- 158
        19851 => X"9D",  -- 157
        19852 => X"9B",  -- 155
        19853 => X"9B",  -- 155
        19854 => X"9D",  -- 157
        19855 => X"9D",  -- 157
        19856 => X"9C",  -- 156
        19857 => X"A5",  -- 165
        19858 => X"A2",  -- 162
        19859 => X"75",  -- 117
        19860 => X"39",  -- 57
        19861 => X"50",  -- 80
        19862 => X"5A",  -- 90
        19863 => X"50",  -- 80
        19864 => X"50",  -- 80
        19865 => X"4B",  -- 75
        19866 => X"43",  -- 67
        19867 => X"3A",  -- 58
        19868 => X"36",  -- 54
        19869 => X"34",  -- 52
        19870 => X"37",  -- 55
        19871 => X"3A",  -- 58
        19872 => X"27",  -- 39
        19873 => X"48",  -- 72
        19874 => X"35",  -- 53
        19875 => X"46",  -- 70
        19876 => X"2A",  -- 42
        19877 => X"3F",  -- 63
        19878 => X"19",  -- 25
        19879 => X"19",  -- 25
        19880 => X"20",  -- 32
        19881 => X"2D",  -- 45
        19882 => X"2B",  -- 43
        19883 => X"2B",  -- 43
        19884 => X"37",  -- 55
        19885 => X"2D",  -- 45
        19886 => X"27",  -- 39
        19887 => X"3B",  -- 59
        19888 => X"4D",  -- 77
        19889 => X"54",  -- 84
        19890 => X"60",  -- 96
        19891 => X"69",  -- 105
        19892 => X"5A",  -- 90
        19893 => X"4F",  -- 79
        19894 => X"5F",  -- 95
        19895 => X"5B",  -- 91
        19896 => X"42",  -- 66
        19897 => X"39",  -- 57
        19898 => X"2D",  -- 45
        19899 => X"4E",  -- 78
        19900 => X"62",  -- 98
        19901 => X"52",  -- 82
        19902 => X"71",  -- 113
        19903 => X"85",  -- 133
        19904 => X"B0",  -- 176
        19905 => X"A4",  -- 164
        19906 => X"97",  -- 151
        19907 => X"87",  -- 135
        19908 => X"6F",  -- 111
        19909 => X"70",  -- 112
        19910 => X"65",  -- 101
        19911 => X"82",  -- 130
        19912 => X"88",  -- 136
        19913 => X"95",  -- 149
        19914 => X"A1",  -- 161
        19915 => X"97",  -- 151
        19916 => X"75",  -- 117
        19917 => X"45",  -- 69
        19918 => X"1F",  -- 31
        19919 => X"0D",  -- 13
        19920 => X"12",  -- 18
        19921 => X"1E",  -- 30
        19922 => X"23",  -- 35
        19923 => X"1D",  -- 29
        19924 => X"15",  -- 21
        19925 => X"15",  -- 21
        19926 => X"15",  -- 21
        19927 => X"14",  -- 20
        19928 => X"11",  -- 17
        19929 => X"08",  -- 8
        19930 => X"10",  -- 16
        19931 => X"21",  -- 33
        19932 => X"40",  -- 64
        19933 => X"5D",  -- 93
        19934 => X"53",  -- 83
        19935 => X"3F",  -- 63
        19936 => X"32",  -- 50
        19937 => X"66",  -- 102
        19938 => X"61",  -- 97
        19939 => X"84",  -- 132
        19940 => X"92",  -- 146
        19941 => X"87",  -- 135
        19942 => X"81",  -- 129
        19943 => X"87",  -- 135
        19944 => X"91",  -- 145
        19945 => X"6D",  -- 109
        19946 => X"3E",  -- 62
        19947 => X"1F",  -- 31
        19948 => X"11",  -- 17
        19949 => X"0A",  -- 10
        19950 => X"0B",  -- 11
        19951 => X"0F",  -- 15
        19952 => X"0C",  -- 12
        19953 => X"0D",  -- 13
        19954 => X"0B",  -- 11
        19955 => X"0E",  -- 14
        19956 => X"1D",  -- 29
        19957 => X"35",  -- 53
        19958 => X"62",  -- 98
        19959 => X"90",  -- 144
        19960 => X"8D",  -- 141
        19961 => X"A9",  -- 169
        19962 => X"B1",  -- 177
        19963 => X"A6",  -- 166
        19964 => X"A6",  -- 166
        19965 => X"B0",  -- 176
        19966 => X"B0",  -- 176
        19967 => X"AD",  -- 173
        19968 => X"A5",  -- 165
        19969 => X"8F",  -- 143
        19970 => X"6C",  -- 108
        19971 => X"45",  -- 69
        19972 => X"49",  -- 73
        19973 => X"25",  -- 37
        19974 => X"1B",  -- 27
        19975 => X"20",  -- 32
        19976 => X"24",  -- 36
        19977 => X"3C",  -- 60
        19978 => X"3E",  -- 62
        19979 => X"34",  -- 52
        19980 => X"54",  -- 84
        19981 => X"4F",  -- 79
        19982 => X"4C",  -- 76
        19983 => X"56",  -- 86
        19984 => X"44",  -- 68
        19985 => X"26",  -- 38
        19986 => X"12",  -- 18
        19987 => X"25",  -- 37
        19988 => X"35",  -- 53
        19989 => X"3C",  -- 60
        19990 => X"38",  -- 56
        19991 => X"3B",  -- 59
        19992 => X"6E",  -- 110
        19993 => X"5F",  -- 95
        19994 => X"77",  -- 119
        19995 => X"81",  -- 129
        19996 => X"44",  -- 68
        19997 => X"3F",  -- 63
        19998 => X"71",  -- 113
        19999 => X"3B",  -- 59
        20000 => X"3A",  -- 58
        20001 => X"36",  -- 54
        20002 => X"47",  -- 71
        20003 => X"3B",  -- 59
        20004 => X"2B",  -- 43
        20005 => X"38",  -- 56
        20006 => X"40",  -- 64
        20007 => X"53",  -- 83
        20008 => X"54",  -- 84
        20009 => X"5E",  -- 94
        20010 => X"49",  -- 73
        20011 => X"31",  -- 49
        20012 => X"55",  -- 85
        20013 => X"BE",  -- 190
        20014 => X"C3",  -- 195
        20015 => X"C1",  -- 193
        20016 => X"B5",  -- 181
        20017 => X"A5",  -- 165
        20018 => X"91",  -- 145
        20019 => X"84",  -- 132
        20020 => X"80",  -- 128
        20021 => X"7E",  -- 126
        20022 => X"79",  -- 121
        20023 => X"73",  -- 115
        20024 => X"78",  -- 120
        20025 => X"76",  -- 118
        20026 => X"78",  -- 120
        20027 => X"7D",  -- 125
        20028 => X"83",  -- 131
        20029 => X"89",  -- 137
        20030 => X"88",  -- 136
        20031 => X"88",  -- 136
        20032 => X"87",  -- 135
        20033 => X"8C",  -- 140
        20034 => X"94",  -- 148
        20035 => X"93",  -- 147
        20036 => X"8A",  -- 138
        20037 => X"82",  -- 130
        20038 => X"88",  -- 136
        20039 => X"93",  -- 147
        20040 => X"99",  -- 153
        20041 => X"A1",  -- 161
        20042 => X"A8",  -- 168
        20043 => X"A8",  -- 168
        20044 => X"A3",  -- 163
        20045 => X"A2",  -- 162
        20046 => X"AA",  -- 170
        20047 => X"B2",  -- 178
        20048 => X"B8",  -- 184
        20049 => X"BB",  -- 187
        20050 => X"BB",  -- 187
        20051 => X"B9",  -- 185
        20052 => X"B4",  -- 180
        20053 => X"B1",  -- 177
        20054 => X"B2",  -- 178
        20055 => X"B4",  -- 180
        20056 => X"B7",  -- 183
        20057 => X"B7",  -- 183
        20058 => X"B3",  -- 179
        20059 => X"A5",  -- 165
        20060 => X"8D",  -- 141
        20061 => X"79",  -- 121
        20062 => X"7C",  -- 124
        20063 => X"88",  -- 136
        20064 => X"A8",  -- 168
        20065 => X"AC",  -- 172
        20066 => X"B2",  -- 178
        20067 => X"B4",  -- 180
        20068 => X"B2",  -- 178
        20069 => X"B0",  -- 176
        20070 => X"AD",  -- 173
        20071 => X"AD",  -- 173
        20072 => X"A8",  -- 168
        20073 => X"A7",  -- 167
        20074 => X"A3",  -- 163
        20075 => X"9E",  -- 158
        20076 => X"9A",  -- 154
        20077 => X"99",  -- 153
        20078 => X"95",  -- 149
        20079 => X"91",  -- 145
        20080 => X"86",  -- 134
        20081 => X"89",  -- 137
        20082 => X"8D",  -- 141
        20083 => X"90",  -- 144
        20084 => X"8A",  -- 138
        20085 => X"73",  -- 115
        20086 => X"4F",  -- 79
        20087 => X"33",  -- 51
        20088 => X"29",  -- 41
        20089 => X"33",  -- 51
        20090 => X"4A",  -- 74
        20091 => X"69",  -- 105
        20092 => X"88",  -- 136
        20093 => X"9D",  -- 157
        20094 => X"A2",  -- 162
        20095 => X"A1",  -- 161
        20096 => X"92",  -- 146
        20097 => X"94",  -- 148
        20098 => X"94",  -- 148
        20099 => X"94",  -- 148
        20100 => X"93",  -- 147
        20101 => X"95",  -- 149
        20102 => X"9C",  -- 156
        20103 => X"A1",  -- 161
        20104 => X"A7",  -- 167
        20105 => X"A8",  -- 168
        20106 => X"A5",  -- 165
        20107 => X"A2",  -- 162
        20108 => X"A1",  -- 161
        20109 => X"A6",  -- 166
        20110 => X"A7",  -- 167
        20111 => X"A5",  -- 165
        20112 => X"9D",  -- 157
        20113 => X"99",  -- 153
        20114 => X"90",  -- 144
        20115 => X"7B",  -- 123
        20116 => X"57",  -- 87
        20117 => X"2F",  -- 47
        20118 => X"1D",  -- 29
        20119 => X"1C",  -- 28
        20120 => X"2C",  -- 44
        20121 => X"48",  -- 72
        20122 => X"67",  -- 103
        20123 => X"79",  -- 121
        20124 => X"81",  -- 129
        20125 => X"86",  -- 134
        20126 => X"8B",  -- 139
        20127 => X"8C",  -- 140
        20128 => X"85",  -- 133
        20129 => X"89",  -- 137
        20130 => X"8A",  -- 138
        20131 => X"85",  -- 133
        20132 => X"7A",  -- 122
        20133 => X"68",  -- 104
        20134 => X"69",  -- 105
        20135 => X"7E",  -- 126
        20136 => X"93",  -- 147
        20137 => X"A3",  -- 163
        20138 => X"A7",  -- 167
        20139 => X"A7",  -- 167
        20140 => X"AC",  -- 172
        20141 => X"AA",  -- 170
        20142 => X"9C",  -- 156
        20143 => X"95",  -- 149
        20144 => X"8B",  -- 139
        20145 => X"8C",  -- 140
        20146 => X"93",  -- 147
        20147 => X"A2",  -- 162
        20148 => X"B2",  -- 178
        20149 => X"B7",  -- 183
        20150 => X"B4",  -- 180
        20151 => X"AF",  -- 175
        20152 => X"AB",  -- 171
        20153 => X"BA",  -- 186
        20154 => X"C1",  -- 193
        20155 => X"BF",  -- 191
        20156 => X"BE",  -- 190
        20157 => X"B6",  -- 182
        20158 => X"AA",  -- 170
        20159 => X"A7",  -- 167
        20160 => X"AB",  -- 171
        20161 => X"AA",  -- 170
        20162 => X"A9",  -- 169
        20163 => X"A9",  -- 169
        20164 => X"A9",  -- 169
        20165 => X"AA",  -- 170
        20166 => X"AA",  -- 170
        20167 => X"A9",  -- 169
        20168 => X"A8",  -- 168
        20169 => X"A6",  -- 166
        20170 => X"A2",  -- 162
        20171 => X"A0",  -- 160
        20172 => X"A0",  -- 160
        20173 => X"A0",  -- 160
        20174 => X"A2",  -- 162
        20175 => X"A3",  -- 163
        20176 => X"AA",  -- 170
        20177 => X"9B",  -- 155
        20178 => X"A6",  -- 166
        20179 => X"A6",  -- 166
        20180 => X"64",  -- 100
        20181 => X"3D",  -- 61
        20182 => X"54",  -- 84
        20183 => X"50",  -- 80
        20184 => X"53",  -- 83
        20185 => X"50",  -- 80
        20186 => X"4A",  -- 74
        20187 => X"40",  -- 64
        20188 => X"36",  -- 54
        20189 => X"2E",  -- 46
        20190 => X"2E",  -- 46
        20191 => X"30",  -- 48
        20192 => X"2D",  -- 45
        20193 => X"28",  -- 40
        20194 => X"3B",  -- 59
        20195 => X"30",  -- 48
        20196 => X"28",  -- 40
        20197 => X"14",  -- 20
        20198 => X"20",  -- 32
        20199 => X"1E",  -- 30
        20200 => X"33",  -- 51
        20201 => X"36",  -- 54
        20202 => X"2A",  -- 42
        20203 => X"33",  -- 51
        20204 => X"4F",  -- 79
        20205 => X"4F",  -- 79
        20206 => X"4D",  -- 77
        20207 => X"66",  -- 102
        20208 => X"8B",  -- 139
        20209 => X"90",  -- 144
        20210 => X"8A",  -- 138
        20211 => X"7C",  -- 124
        20212 => X"65",  -- 101
        20213 => X"62",  -- 98
        20214 => X"67",  -- 103
        20215 => X"4E",  -- 78
        20216 => X"46",  -- 70
        20217 => X"3A",  -- 58
        20218 => X"28",  -- 40
        20219 => X"69",  -- 105
        20220 => X"78",  -- 120
        20221 => X"7A",  -- 122
        20222 => X"87",  -- 135
        20223 => X"66",  -- 102
        20224 => X"67",  -- 103
        20225 => X"74",  -- 116
        20226 => X"76",  -- 118
        20227 => X"6F",  -- 111
        20228 => X"68",  -- 104
        20229 => X"7A",  -- 122
        20230 => X"6B",  -- 107
        20231 => X"87",  -- 135
        20232 => X"9B",  -- 155
        20233 => X"91",  -- 145
        20234 => X"79",  -- 121
        20235 => X"5A",  -- 90
        20236 => X"33",  -- 51
        20237 => X"1C",  -- 28
        20238 => X"12",  -- 18
        20239 => X"16",  -- 22
        20240 => X"20",  -- 32
        20241 => X"2B",  -- 43
        20242 => X"2D",  -- 45
        20243 => X"1F",  -- 31
        20244 => X"14",  -- 20
        20245 => X"13",  -- 19
        20246 => X"0E",  -- 14
        20247 => X"05",  -- 5
        20248 => X"0C",  -- 12
        20249 => X"0D",  -- 13
        20250 => X"17",  -- 23
        20251 => X"2A",  -- 42
        20252 => X"3F",  -- 63
        20253 => X"51",  -- 81
        20254 => X"56",  -- 86
        20255 => X"48",  -- 72
        20256 => X"38",  -- 56
        20257 => X"7A",  -- 122
        20258 => X"67",  -- 103
        20259 => X"75",  -- 117
        20260 => X"8A",  -- 138
        20261 => X"8A",  -- 138
        20262 => X"89",  -- 137
        20263 => X"8C",  -- 140
        20264 => X"79",  -- 121
        20265 => X"8C",  -- 140
        20266 => X"60",  -- 96
        20267 => X"26",  -- 38
        20268 => X"1D",  -- 29
        20269 => X"16",  -- 22
        20270 => X"06",  -- 6
        20271 => X"0E",  -- 14
        20272 => X"12",  -- 18
        20273 => X"0E",  -- 14
        20274 => X"09",  -- 9
        20275 => X"0C",  -- 12
        20276 => X"15",  -- 21
        20277 => X"1D",  -- 29
        20278 => X"34",  -- 52
        20279 => X"53",  -- 83
        20280 => X"89",  -- 137
        20281 => X"90",  -- 144
        20282 => X"8E",  -- 142
        20283 => X"8D",  -- 141
        20284 => X"95",  -- 149
        20285 => X"99",  -- 153
        20286 => X"9E",  -- 158
        20287 => X"A7",  -- 167
        20288 => X"AC",  -- 172
        20289 => X"A0",  -- 160
        20290 => X"72",  -- 114
        20291 => X"4C",  -- 76
        20292 => X"4C",  -- 76
        20293 => X"42",  -- 66
        20294 => X"2C",  -- 44
        20295 => X"2A",  -- 42
        20296 => X"3C",  -- 60
        20297 => X"38",  -- 56
        20298 => X"44",  -- 68
        20299 => X"47",  -- 71
        20300 => X"43",  -- 67
        20301 => X"24",  -- 36
        20302 => X"2C",  -- 44
        20303 => X"42",  -- 66
        20304 => X"2A",  -- 42
        20305 => X"2B",  -- 43
        20306 => X"30",  -- 48
        20307 => X"38",  -- 56
        20308 => X"44",  -- 68
        20309 => X"48",  -- 72
        20310 => X"47",  -- 71
        20311 => X"44",  -- 68
        20312 => X"54",  -- 84
        20313 => X"62",  -- 98
        20314 => X"73",  -- 115
        20315 => X"7B",  -- 123
        20316 => X"5B",  -- 91
        20317 => X"22",  -- 34
        20318 => X"39",  -- 57
        20319 => X"4B",  -- 75
        20320 => X"48",  -- 72
        20321 => X"3F",  -- 63
        20322 => X"31",  -- 49
        20323 => X"37",  -- 55
        20324 => X"35",  -- 53
        20325 => X"39",  -- 57
        20326 => X"46",  -- 70
        20327 => X"44",  -- 68
        20328 => X"48",  -- 72
        20329 => X"3D",  -- 61
        20330 => X"22",  -- 34
        20331 => X"33",  -- 51
        20332 => X"B3",  -- 179
        20333 => X"C2",  -- 194
        20334 => X"C1",  -- 193
        20335 => X"BD",  -- 189
        20336 => X"B5",  -- 181
        20337 => X"A2",  -- 162
        20338 => X"8A",  -- 138
        20339 => X"7C",  -- 124
        20340 => X"7B",  -- 123
        20341 => X"7C",  -- 124
        20342 => X"79",  -- 121
        20343 => X"75",  -- 117
        20344 => X"77",  -- 119
        20345 => X"74",  -- 116
        20346 => X"72",  -- 114
        20347 => X"73",  -- 115
        20348 => X"7A",  -- 122
        20349 => X"7E",  -- 126
        20350 => X"7F",  -- 127
        20351 => X"7F",  -- 127
        20352 => X"8E",  -- 142
        20353 => X"8B",  -- 139
        20354 => X"8C",  -- 140
        20355 => X"90",  -- 144
        20356 => X"91",  -- 145
        20357 => X"93",  -- 147
        20358 => X"9B",  -- 155
        20359 => X"A5",  -- 165
        20360 => X"AC",  -- 172
        20361 => X"AC",  -- 172
        20362 => X"A9",  -- 169
        20363 => X"A4",  -- 164
        20364 => X"A1",  -- 161
        20365 => X"A1",  -- 161
        20366 => X"A5",  -- 165
        20367 => X"AA",  -- 170
        20368 => X"B1",  -- 177
        20369 => X"B4",  -- 180
        20370 => X"B8",  -- 184
        20371 => X"BA",  -- 186
        20372 => X"BA",  -- 186
        20373 => X"BA",  -- 186
        20374 => X"B8",  -- 184
        20375 => X"B8",  -- 184
        20376 => X"BE",  -- 190
        20377 => X"BA",  -- 186
        20378 => X"BC",  -- 188
        20379 => X"B7",  -- 183
        20380 => X"9B",  -- 155
        20381 => X"7C",  -- 124
        20382 => X"7B",  -- 123
        20383 => X"8D",  -- 141
        20384 => X"A5",  -- 165
        20385 => X"A9",  -- 169
        20386 => X"AE",  -- 174
        20387 => X"B1",  -- 177
        20388 => X"B1",  -- 177
        20389 => X"AF",  -- 175
        20390 => X"AD",  -- 173
        20391 => X"AC",  -- 172
        20392 => X"A6",  -- 166
        20393 => X"AA",  -- 170
        20394 => X"A8",  -- 168
        20395 => X"A2",  -- 162
        20396 => X"A3",  -- 163
        20397 => X"A4",  -- 164
        20398 => X"9C",  -- 156
        20399 => X"91",  -- 145
        20400 => X"8C",  -- 140
        20401 => X"8B",  -- 139
        20402 => X"8D",  -- 141
        20403 => X"8F",  -- 143
        20404 => X"8C",  -- 140
        20405 => X"78",  -- 120
        20406 => X"60",  -- 96
        20407 => X"4E",  -- 78
        20408 => X"2D",  -- 45
        20409 => X"3C",  -- 60
        20410 => X"54",  -- 84
        20411 => X"6E",  -- 110
        20412 => X"83",  -- 131
        20413 => X"91",  -- 145
        20414 => X"9A",  -- 154
        20415 => X"9D",  -- 157
        20416 => X"94",  -- 148
        20417 => X"96",  -- 150
        20418 => X"97",  -- 151
        20419 => X"97",  -- 151
        20420 => X"96",  -- 150
        20421 => X"99",  -- 153
        20422 => X"A0",  -- 160
        20423 => X"A5",  -- 165
        20424 => X"A9",  -- 169
        20425 => X"AB",  -- 171
        20426 => X"A8",  -- 168
        20427 => X"A0",  -- 160
        20428 => X"9F",  -- 159
        20429 => X"A2",  -- 162
        20430 => X"A4",  -- 164
        20431 => X"A4",  -- 164
        20432 => X"9E",  -- 158
        20433 => X"9F",  -- 159
        20434 => X"96",  -- 150
        20435 => X"75",  -- 117
        20436 => X"46",  -- 70
        20437 => X"23",  -- 35
        20438 => X"1C",  -- 28
        20439 => X"22",  -- 34
        20440 => X"36",  -- 54
        20441 => X"4D",  -- 77
        20442 => X"69",  -- 105
        20443 => X"78",  -- 120
        20444 => X"82",  -- 130
        20445 => X"8B",  -- 139
        20446 => X"90",  -- 144
        20447 => X"90",  -- 144
        20448 => X"8A",  -- 138
        20449 => X"8C",  -- 140
        20450 => X"8B",  -- 139
        20451 => X"85",  -- 133
        20452 => X"7C",  -- 124
        20453 => X"6E",  -- 110
        20454 => X"76",  -- 118
        20455 => X"90",  -- 144
        20456 => X"9D",  -- 157
        20457 => X"AC",  -- 172
        20458 => X"AE",  -- 174
        20459 => X"AC",  -- 172
        20460 => X"AD",  -- 173
        20461 => X"A7",  -- 167
        20462 => X"97",  -- 151
        20463 => X"8F",  -- 143
        20464 => X"91",  -- 145
        20465 => X"90",  -- 144
        20466 => X"96",  -- 150
        20467 => X"A3",  -- 163
        20468 => X"B1",  -- 177
        20469 => X"B3",  -- 179
        20470 => X"AB",  -- 171
        20471 => X"A3",  -- 163
        20472 => X"A9",  -- 169
        20473 => X"BC",  -- 188
        20474 => X"C2",  -- 194
        20475 => X"C1",  -- 193
        20476 => X"C1",  -- 193
        20477 => X"BB",  -- 187
        20478 => X"B0",  -- 176
        20479 => X"AF",  -- 175
        20480 => X"AD",  -- 173
        20481 => X"AD",  -- 173
        20482 => X"AF",  -- 175
        20483 => X"AF",  -- 175
        20484 => X"AF",  -- 175
        20485 => X"AE",  -- 174
        20486 => X"AD",  -- 173
        20487 => X"AC",  -- 172
        20488 => X"A8",  -- 168
        20489 => X"A9",  -- 169
        20490 => X"A8",  -- 168
        20491 => X"A5",  -- 165
        20492 => X"A2",  -- 162
        20493 => X"A1",  -- 161
        20494 => X"A2",  -- 162
        20495 => X"A6",  -- 166
        20496 => X"A7",  -- 167
        20497 => X"A3",  -- 163
        20498 => X"A7",  -- 167
        20499 => X"AB",  -- 171
        20500 => X"91",  -- 145
        20501 => X"61",  -- 97
        20502 => X"3E",  -- 62
        20503 => X"35",  -- 53
        20504 => X"3D",  -- 61
        20505 => X"4A",  -- 74
        20506 => X"3F",  -- 63
        20507 => X"33",  -- 51
        20508 => X"39",  -- 57
        20509 => X"31",  -- 49
        20510 => X"26",  -- 38
        20511 => X"34",  -- 52
        20512 => X"30",  -- 48
        20513 => X"34",  -- 52
        20514 => X"40",  -- 64
        20515 => X"3A",  -- 58
        20516 => X"30",  -- 48
        20517 => X"3D",  -- 61
        20518 => X"41",  -- 65
        20519 => X"2C",  -- 44
        20520 => X"38",  -- 56
        20521 => X"4C",  -- 76
        20522 => X"4C",  -- 76
        20523 => X"3D",  -- 61
        20524 => X"44",  -- 68
        20525 => X"57",  -- 87
        20526 => X"63",  -- 99
        20527 => X"68",  -- 104
        20528 => X"5E",  -- 94
        20529 => X"5E",  -- 94
        20530 => X"52",  -- 82
        20531 => X"44",  -- 68
        20532 => X"51",  -- 81
        20533 => X"67",  -- 103
        20534 => X"63",  -- 99
        20535 => X"4C",  -- 76
        20536 => X"35",  -- 53
        20537 => X"43",  -- 67
        20538 => X"6F",  -- 111
        20539 => X"7B",  -- 123
        20540 => X"7B",  -- 123
        20541 => X"74",  -- 116
        20542 => X"6D",  -- 109
        20543 => X"46",  -- 70
        20544 => X"28",  -- 40
        20545 => X"2A",  -- 42
        20546 => X"45",  -- 69
        20547 => X"70",  -- 112
        20548 => X"85",  -- 133
        20549 => X"81",  -- 129
        20550 => X"81",  -- 129
        20551 => X"8C",  -- 140
        20552 => X"96",  -- 150
        20553 => X"81",  -- 129
        20554 => X"40",  -- 64
        20555 => X"30",  -- 48
        20556 => X"12",  -- 18
        20557 => X"0D",  -- 13
        20558 => X"16",  -- 22
        20559 => X"19",  -- 25
        20560 => X"27",  -- 39
        20561 => X"21",  -- 33
        20562 => X"1A",  -- 26
        20563 => X"16",  -- 22
        20564 => X"0D",  -- 13
        20565 => X"08",  -- 8
        20566 => X"0D",  -- 13
        20567 => X"16",  -- 22
        20568 => X"1A",  -- 26
        20569 => X"1B",  -- 27
        20570 => X"55",  -- 85
        20571 => X"64",  -- 100
        20572 => X"63",  -- 99
        20573 => X"65",  -- 101
        20574 => X"5F",  -- 95
        20575 => X"33",  -- 51
        20576 => X"31",  -- 49
        20577 => X"76",  -- 118
        20578 => X"7C",  -- 124
        20579 => X"6A",  -- 106
        20580 => X"70",  -- 112
        20581 => X"91",  -- 145
        20582 => X"85",  -- 133
        20583 => X"86",  -- 134
        20584 => X"82",  -- 130
        20585 => X"87",  -- 135
        20586 => X"87",  -- 135
        20587 => X"62",  -- 98
        20588 => X"51",  -- 81
        20589 => X"34",  -- 52
        20590 => X"25",  -- 37
        20591 => X"0B",  -- 11
        20592 => X"07",  -- 7
        20593 => X"0E",  -- 14
        20594 => X"12",  -- 18
        20595 => X"11",  -- 17
        20596 => X"11",  -- 17
        20597 => X"17",  -- 23
        20598 => X"1B",  -- 27
        20599 => X"1D",  -- 29
        20600 => X"45",  -- 69
        20601 => X"6D",  -- 109
        20602 => X"8A",  -- 138
        20603 => X"8C",  -- 140
        20604 => X"81",  -- 129
        20605 => X"77",  -- 119
        20606 => X"79",  -- 121
        20607 => X"84",  -- 132
        20608 => X"8C",  -- 140
        20609 => X"8A",  -- 138
        20610 => X"6C",  -- 108
        20611 => X"42",  -- 66
        20612 => X"3E",  -- 62
        20613 => X"55",  -- 85
        20614 => X"52",  -- 82
        20615 => X"34",  -- 52
        20616 => X"2E",  -- 46
        20617 => X"3B",  -- 59
        20618 => X"48",  -- 72
        20619 => X"54",  -- 84
        20620 => X"4F",  -- 79
        20621 => X"3D",  -- 61
        20622 => X"40",  -- 64
        20623 => X"57",  -- 87
        20624 => X"5A",  -- 90
        20625 => X"4C",  -- 76
        20626 => X"41",  -- 65
        20627 => X"5A",  -- 90
        20628 => X"70",  -- 112
        20629 => X"6B",  -- 107
        20630 => X"61",  -- 97
        20631 => X"4F",  -- 79
        20632 => X"57",  -- 87
        20633 => X"44",  -- 68
        20634 => X"66",  -- 102
        20635 => X"73",  -- 115
        20636 => X"42",  -- 66
        20637 => X"4F",  -- 79
        20638 => X"26",  -- 38
        20639 => X"4F",  -- 79
        20640 => X"67",  -- 103
        20641 => X"4C",  -- 76
        20642 => X"30",  -- 48
        20643 => X"30",  -- 48
        20644 => X"35",  -- 53
        20645 => X"37",  -- 55
        20646 => X"40",  -- 64
        20647 => X"35",  -- 53
        20648 => X"25",  -- 37
        20649 => X"0F",  -- 15
        20650 => X"49",  -- 73
        20651 => X"B2",  -- 178
        20652 => X"D3",  -- 211
        20653 => X"BA",  -- 186
        20654 => X"BC",  -- 188
        20655 => X"CE",  -- 206
        20656 => X"C4",  -- 196
        20657 => X"A8",  -- 168
        20658 => X"8C",  -- 140
        20659 => X"83",  -- 131
        20660 => X"8C",  -- 140
        20661 => X"8F",  -- 143
        20662 => X"80",  -- 128
        20663 => X"6C",  -- 108
        20664 => X"7D",  -- 125
        20665 => X"7A",  -- 122
        20666 => X"77",  -- 119
        20667 => X"79",  -- 121
        20668 => X"80",  -- 128
        20669 => X"84",  -- 132
        20670 => X"84",  -- 132
        20671 => X"81",  -- 129
        20672 => X"81",  -- 129
        20673 => X"89",  -- 137
        20674 => X"93",  -- 147
        20675 => X"97",  -- 151
        20676 => X"98",  -- 152
        20677 => X"98",  -- 152
        20678 => X"9B",  -- 155
        20679 => X"9F",  -- 159
        20680 => X"A3",  -- 163
        20681 => X"A1",  -- 161
        20682 => X"A2",  -- 162
        20683 => X"A5",  -- 165
        20684 => X"A6",  -- 166
        20685 => X"A8",  -- 168
        20686 => X"AF",  -- 175
        20687 => X"B6",  -- 182
        20688 => X"BB",  -- 187
        20689 => X"BB",  -- 187
        20690 => X"BD",  -- 189
        20691 => X"BE",  -- 190
        20692 => X"BF",  -- 191
        20693 => X"C1",  -- 193
        20694 => X"C5",  -- 197
        20695 => X"C7",  -- 199
        20696 => X"BE",  -- 190
        20697 => X"BE",  -- 190
        20698 => X"B9",  -- 185
        20699 => X"A9",  -- 169
        20700 => X"8E",  -- 142
        20701 => X"7D",  -- 125
        20702 => X"80",  -- 128
        20703 => X"8E",  -- 142
        20704 => X"96",  -- 150
        20705 => X"A5",  -- 165
        20706 => X"B3",  -- 179
        20707 => X"B8",  -- 184
        20708 => X"B7",  -- 183
        20709 => X"B4",  -- 180
        20710 => X"AE",  -- 174
        20711 => X"A9",  -- 169
        20712 => X"AA",  -- 170
        20713 => X"A6",  -- 166
        20714 => X"A2",  -- 162
        20715 => X"A1",  -- 161
        20716 => X"A3",  -- 163
        20717 => X"A3",  -- 163
        20718 => X"9F",  -- 159
        20719 => X"9B",  -- 155
        20720 => X"9A",  -- 154
        20721 => X"91",  -- 145
        20722 => X"8E",  -- 142
        20723 => X"90",  -- 144
        20724 => X"8B",  -- 139
        20725 => X"7E",  -- 126
        20726 => X"62",  -- 98
        20727 => X"40",  -- 64
        20728 => X"25",  -- 37
        20729 => X"3B",  -- 59
        20730 => X"5E",  -- 94
        20731 => X"74",  -- 116
        20732 => X"7A",  -- 122
        20733 => X"7C",  -- 124
        20734 => X"89",  -- 137
        20735 => X"98",  -- 152
        20736 => X"9C",  -- 156
        20737 => X"98",  -- 152
        20738 => X"92",  -- 146
        20739 => X"90",  -- 144
        20740 => X"90",  -- 144
        20741 => X"96",  -- 150
        20742 => X"9B",  -- 155
        20743 => X"A1",  -- 161
        20744 => X"99",  -- 153
        20745 => X"97",  -- 151
        20746 => X"99",  -- 153
        20747 => X"9E",  -- 158
        20748 => X"A7",  -- 167
        20749 => X"AA",  -- 170
        20750 => X"A5",  -- 165
        20751 => X"A1",  -- 161
        20752 => X"A9",  -- 169
        20753 => X"9F",  -- 159
        20754 => X"92",  -- 146
        20755 => X"7D",  -- 125
        20756 => X"59",  -- 89
        20757 => X"33",  -- 51
        20758 => X"26",  -- 38
        20759 => X"2D",  -- 45
        20760 => X"32",  -- 50
        20761 => X"50",  -- 80
        20762 => X"70",  -- 112
        20763 => X"84",  -- 132
        20764 => X"8D",  -- 141
        20765 => X"90",  -- 144
        20766 => X"8E",  -- 142
        20767 => X"88",  -- 136
        20768 => X"81",  -- 129
        20769 => X"8E",  -- 142
        20770 => X"94",  -- 148
        20771 => X"89",  -- 137
        20772 => X"79",  -- 121
        20773 => X"75",  -- 117
        20774 => X"81",  -- 129
        20775 => X"8E",  -- 142
        20776 => X"9C",  -- 156
        20777 => X"9E",  -- 158
        20778 => X"A6",  -- 166
        20779 => X"AC",  -- 172
        20780 => X"A9",  -- 169
        20781 => X"9E",  -- 158
        20782 => X"92",  -- 146
        20783 => X"8D",  -- 141
        20784 => X"9A",  -- 154
        20785 => X"9B",  -- 155
        20786 => X"A2",  -- 162
        20787 => X"AE",  -- 174
        20788 => X"B3",  -- 179
        20789 => X"A9",  -- 169
        20790 => X"97",  -- 151
        20791 => X"89",  -- 137
        20792 => X"9E",  -- 158
        20793 => X"B7",  -- 183
        20794 => X"C6",  -- 198
        20795 => X"C3",  -- 195
        20796 => X"C0",  -- 192
        20797 => X"B9",  -- 185
        20798 => X"B5",  -- 181
        20799 => X"B8",  -- 184
        20800 => X"AB",  -- 171
        20801 => X"AE",  -- 174
        20802 => X"B0",  -- 176
        20803 => X"B3",  -- 179
        20804 => X"B3",  -- 179
        20805 => X"B2",  -- 178
        20806 => X"AE",  -- 174
        20807 => X"AC",  -- 172
        20808 => X"A9",  -- 169
        20809 => X"AA",  -- 170
        20810 => X"AA",  -- 170
        20811 => X"A8",  -- 168
        20812 => X"A6",  -- 166
        20813 => X"A4",  -- 164
        20814 => X"A6",  -- 166
        20815 => X"A8",  -- 168
        20816 => X"A6",  -- 166
        20817 => X"AA",  -- 170
        20818 => X"A7",  -- 167
        20819 => X"A2",  -- 162
        20820 => X"A3",  -- 163
        20821 => X"93",  -- 147
        20822 => X"5E",  -- 94
        20823 => X"26",  -- 38
        20824 => X"2E",  -- 46
        20825 => X"3A",  -- 58
        20826 => X"38",  -- 56
        20827 => X"34",  -- 52
        20828 => X"3A",  -- 58
        20829 => X"33",  -- 51
        20830 => X"27",  -- 39
        20831 => X"2C",  -- 44
        20832 => X"39",  -- 57
        20833 => X"39",  -- 57
        20834 => X"42",  -- 66
        20835 => X"43",  -- 67
        20836 => X"3C",  -- 60
        20837 => X"4D",  -- 77
        20838 => X"62",  -- 98
        20839 => X"65",  -- 101
        20840 => X"6D",  -- 109
        20841 => X"70",  -- 112
        20842 => X"6A",  -- 106
        20843 => X"6A",  -- 106
        20844 => X"6F",  -- 111
        20845 => X"6B",  -- 107
        20846 => X"61",  -- 97
        20847 => X"5E",  -- 94
        20848 => X"45",  -- 69
        20849 => X"51",  -- 81
        20850 => X"56",  -- 86
        20851 => X"4E",  -- 78
        20852 => X"4B",  -- 75
        20853 => X"4B",  -- 75
        20854 => X"45",  -- 69
        20855 => X"38",  -- 56
        20856 => X"3F",  -- 63
        20857 => X"5E",  -- 94
        20858 => X"89",  -- 137
        20859 => X"8E",  -- 142
        20860 => X"89",  -- 137
        20861 => X"5A",  -- 90
        20862 => X"36",  -- 54
        20863 => X"1D",  -- 29
        20864 => X"05",  -- 5
        20865 => X"21",  -- 33
        20866 => X"4E",  -- 78
        20867 => X"73",  -- 115
        20868 => X"82",  -- 130
        20869 => X"83",  -- 131
        20870 => X"87",  -- 135
        20871 => X"8C",  -- 140
        20872 => X"5A",  -- 90
        20873 => X"3F",  -- 63
        20874 => X"1F",  -- 31
        20875 => X"17",  -- 23
        20876 => X"0D",  -- 13
        20877 => X"1A",  -- 26
        20878 => X"12",  -- 18
        20879 => X"18",  -- 24
        20880 => X"1B",  -- 27
        20881 => X"18",  -- 24
        20882 => X"13",  -- 19
        20883 => X"0D",  -- 13
        20884 => X"0A",  -- 10
        20885 => X"13",  -- 19
        20886 => X"26",  -- 38
        20887 => X"38",  -- 56
        20888 => X"4A",  -- 74
        20889 => X"5F",  -- 95
        20890 => X"7B",  -- 123
        20891 => X"82",  -- 130
        20892 => X"6C",  -- 108
        20893 => X"5E",  -- 94
        20894 => X"5D",  -- 93
        20895 => X"2B",  -- 43
        20896 => X"27",  -- 39
        20897 => X"65",  -- 101
        20898 => X"7A",  -- 122
        20899 => X"75",  -- 117
        20900 => X"6E",  -- 110
        20901 => X"7C",  -- 124
        20902 => X"78",  -- 120
        20903 => X"83",  -- 131
        20904 => X"84",  -- 132
        20905 => X"8A",  -- 138
        20906 => X"96",  -- 150
        20907 => X"89",  -- 137
        20908 => X"89",  -- 137
        20909 => X"72",  -- 114
        20910 => X"5E",  -- 94
        20911 => X"43",  -- 67
        20912 => X"26",  -- 38
        20913 => X"18",  -- 24
        20914 => X"0F",  -- 15
        20915 => X"10",  -- 16
        20916 => X"10",  -- 16
        20917 => X"0D",  -- 13
        20918 => X"0C",  -- 12
        20919 => X"0F",  -- 15
        20920 => X"1A",  -- 26
        20921 => X"3E",  -- 62
        20922 => X"69",  -- 105
        20923 => X"85",  -- 133
        20924 => X"88",  -- 136
        20925 => X"74",  -- 116
        20926 => X"60",  -- 96
        20927 => X"58",  -- 88
        20928 => X"5D",  -- 93
        20929 => X"54",  -- 84
        20930 => X"3D",  -- 61
        20931 => X"28",  -- 40
        20932 => X"2D",  -- 45
        20933 => X"49",  -- 73
        20934 => X"65",  -- 101
        20935 => X"70",  -- 112
        20936 => X"2B",  -- 43
        20937 => X"26",  -- 38
        20938 => X"3D",  -- 61
        20939 => X"4A",  -- 74
        20940 => X"49",  -- 73
        20941 => X"40",  -- 64
        20942 => X"40",  -- 64
        20943 => X"72",  -- 114
        20944 => X"74",  -- 116
        20945 => X"76",  -- 118
        20946 => X"65",  -- 101
        20947 => X"5B",  -- 91
        20948 => X"5F",  -- 95
        20949 => X"6C",  -- 108
        20950 => X"82",  -- 130
        20951 => X"80",  -- 128
        20952 => X"80",  -- 128
        20953 => X"64",  -- 100
        20954 => X"60",  -- 96
        20955 => X"53",  -- 83
        20956 => X"39",  -- 57
        20957 => X"53",  -- 83
        20958 => X"3E",  -- 62
        20959 => X"59",  -- 89
        20960 => X"5E",  -- 94
        20961 => X"4E",  -- 78
        20962 => X"3A",  -- 58
        20963 => X"2D",  -- 45
        20964 => X"36",  -- 54
        20965 => X"3E",  -- 62
        20966 => X"30",  -- 48
        20967 => X"1F",  -- 31
        20968 => X"16",  -- 22
        20969 => X"66",  -- 102
        20970 => X"A8",  -- 168
        20971 => X"BA",  -- 186
        20972 => X"BF",  -- 191
        20973 => X"CC",  -- 204
        20974 => X"CB",  -- 203
        20975 => X"BF",  -- 191
        20976 => X"B3",  -- 179
        20977 => X"B1",  -- 177
        20978 => X"AB",  -- 171
        20979 => X"A2",  -- 162
        20980 => X"97",  -- 151
        20981 => X"8D",  -- 141
        20982 => X"81",  -- 129
        20983 => X"7C",  -- 124
        20984 => X"7B",  -- 123
        20985 => X"7B",  -- 123
        20986 => X"7E",  -- 126
        20987 => X"86",  -- 134
        20988 => X"8E",  -- 142
        20989 => X"91",  -- 145
        20990 => X"8D",  -- 141
        20991 => X"87",  -- 135
        20992 => X"7B",  -- 123
        20993 => X"7D",  -- 125
        20994 => X"83",  -- 131
        20995 => X"88",  -- 136
        20996 => X"8E",  -- 142
        20997 => X"95",  -- 149
        20998 => X"99",  -- 153
        20999 => X"9A",  -- 154
        21000 => X"9A",  -- 154
        21001 => X"9D",  -- 157
        21002 => X"A1",  -- 161
        21003 => X"A3",  -- 163
        21004 => X"A1",  -- 161
        21005 => X"A2",  -- 162
        21006 => X"AB",  -- 171
        21007 => X"B5",  -- 181
        21008 => X"B6",  -- 182
        21009 => X"BA",  -- 186
        21010 => X"C0",  -- 192
        21011 => X"C4",  -- 196
        21012 => X"C6",  -- 198
        21013 => X"C4",  -- 196
        21014 => X"C4",  -- 196
        21015 => X"C4",  -- 196
        21016 => X"CA",  -- 202
        21017 => X"C8",  -- 200
        21018 => X"C5",  -- 197
        21019 => X"BA",  -- 186
        21020 => X"A8",  -- 168
        21021 => X"95",  -- 149
        21022 => X"8E",  -- 142
        21023 => X"91",  -- 145
        21024 => X"97",  -- 151
        21025 => X"A7",  -- 167
        21026 => X"B6",  -- 182
        21027 => X"BA",  -- 186
        21028 => X"B4",  -- 180
        21029 => X"AF",  -- 175
        21030 => X"AD",  -- 173
        21031 => X"AC",  -- 172
        21032 => X"A8",  -- 168
        21033 => X"A6",  -- 166
        21034 => X"A3",  -- 163
        21035 => X"A4",  -- 164
        21036 => X"A6",  -- 166
        21037 => X"A6",  -- 166
        21038 => X"A2",  -- 162
        21039 => X"A0",  -- 160
        21040 => X"A2",  -- 162
        21041 => X"93",  -- 147
        21042 => X"8B",  -- 139
        21043 => X"86",  -- 134
        21044 => X"7F",  -- 127
        21045 => X"73",  -- 115
        21046 => X"57",  -- 87
        21047 => X"37",  -- 55
        21048 => X"35",  -- 53
        21049 => X"3C",  -- 60
        21050 => X"4F",  -- 79
        21051 => X"6C",  -- 108
        21052 => X"83",  -- 131
        21053 => X"8E",  -- 142
        21054 => X"92",  -- 146
        21055 => X"93",  -- 147
        21056 => X"91",  -- 145
        21057 => X"93",  -- 147
        21058 => X"93",  -- 147
        21059 => X"98",  -- 152
        21060 => X"9B",  -- 155
        21061 => X"9D",  -- 157
        21062 => X"9B",  -- 155
        21063 => X"9A",  -- 154
        21064 => X"9F",  -- 159
        21065 => X"9E",  -- 158
        21066 => X"A0",  -- 160
        21067 => X"A6",  -- 166
        21068 => X"AD",  -- 173
        21069 => X"AF",  -- 175
        21070 => X"AD",  -- 173
        21071 => X"AC",  -- 172
        21072 => X"9D",  -- 157
        21073 => X"A7",  -- 167
        21074 => X"9A",  -- 154
        21075 => X"6B",  -- 107
        21076 => X"37",  -- 55
        21077 => X"1F",  -- 31
        21078 => X"24",  -- 36
        21079 => X"30",  -- 48
        21080 => X"3D",  -- 61
        21081 => X"56",  -- 86
        21082 => X"72",  -- 114
        21083 => X"80",  -- 128
        21084 => X"86",  -- 134
        21085 => X"8D",  -- 141
        21086 => X"92",  -- 146
        21087 => X"90",  -- 144
        21088 => X"8C",  -- 140
        21089 => X"8F",  -- 143
        21090 => X"8B",  -- 139
        21091 => X"7E",  -- 126
        21092 => X"72",  -- 114
        21093 => X"78",  -- 120
        21094 => X"8E",  -- 142
        21095 => X"A4",  -- 164
        21096 => X"A1",  -- 161
        21097 => X"A4",  -- 164
        21098 => X"AB",  -- 171
        21099 => X"AF",  -- 175
        21100 => X"AA",  -- 170
        21101 => X"A0",  -- 160
        21102 => X"9B",  -- 155
        21103 => X"9B",  -- 155
        21104 => X"A3",  -- 163
        21105 => X"A5",  -- 165
        21106 => X"AC",  -- 172
        21107 => X"B3",  -- 179
        21108 => X"B5",  -- 181
        21109 => X"A9",  -- 169
        21110 => X"95",  -- 149
        21111 => X"85",  -- 133
        21112 => X"9B",  -- 155
        21113 => X"B7",  -- 183
        21114 => X"C3",  -- 195
        21115 => X"BC",  -- 188
        21116 => X"B8",  -- 184
        21117 => X"B8",  -- 184
        21118 => X"B8",  -- 184
        21119 => X"BC",  -- 188
        21120 => X"A9",  -- 169
        21121 => X"AC",  -- 172
        21122 => X"AF",  -- 175
        21123 => X"B3",  -- 179
        21124 => X"B3",  -- 179
        21125 => X"AF",  -- 175
        21126 => X"AB",  -- 171
        21127 => X"A9",  -- 169
        21128 => X"A7",  -- 167
        21129 => X"A8",  -- 168
        21130 => X"AA",  -- 170
        21131 => X"A9",  -- 169
        21132 => X"A8",  -- 168
        21133 => X"A7",  -- 167
        21134 => X"A7",  -- 167
        21135 => X"A8",  -- 168
        21136 => X"A2",  -- 162
        21137 => X"AF",  -- 175
        21138 => X"AB",  -- 171
        21139 => X"9D",  -- 157
        21140 => X"A0",  -- 160
        21141 => X"A8",  -- 168
        21142 => X"8C",  -- 140
        21143 => X"5E",  -- 94
        21144 => X"1D",  -- 29
        21145 => X"23",  -- 35
        21146 => X"29",  -- 41
        21147 => X"2D",  -- 45
        21148 => X"30",  -- 48
        21149 => X"32",  -- 50
        21150 => X"35",  -- 53
        21151 => X"3B",  -- 59
        21152 => X"3E",  -- 62
        21153 => X"45",  -- 69
        21154 => X"56",  -- 86
        21155 => X"5D",  -- 93
        21156 => X"50",  -- 80
        21157 => X"4B",  -- 75
        21158 => X"50",  -- 80
        21159 => X"53",  -- 83
        21160 => X"70",  -- 112
        21161 => X"61",  -- 97
        21162 => X"53",  -- 83
        21163 => X"56",  -- 86
        21164 => X"58",  -- 88
        21165 => X"4B",  -- 75
        21166 => X"40",  -- 64
        21167 => X"47",  -- 71
        21168 => X"46",  -- 70
        21169 => X"5B",  -- 91
        21170 => X"5E",  -- 94
        21171 => X"49",  -- 73
        21172 => X"3F",  -- 63
        21173 => X"4B",  -- 75
        21174 => X"52",  -- 82
        21175 => X"4C",  -- 76
        21176 => X"64",  -- 100
        21177 => X"7F",  -- 127
        21178 => X"8E",  -- 142
        21179 => X"78",  -- 120
        21180 => X"67",  -- 103
        21181 => X"29",  -- 41
        21182 => X"0B",  -- 11
        21183 => X"0E",  -- 14
        21184 => X"1F",  -- 31
        21185 => X"37",  -- 55
        21186 => X"56",  -- 86
        21187 => X"73",  -- 115
        21188 => X"89",  -- 137
        21189 => X"8C",  -- 140
        21190 => X"78",  -- 120
        21191 => X"5E",  -- 94
        21192 => X"2F",  -- 47
        21193 => X"15",  -- 21
        21194 => X"0E",  -- 14
        21195 => X"0A",  -- 10
        21196 => X"0F",  -- 15
        21197 => X"26",  -- 38
        21198 => X"0F",  -- 15
        21199 => X"14",  -- 20
        21200 => X"0A",  -- 10
        21201 => X"11",  -- 17
        21202 => X"15",  -- 21
        21203 => X"16",  -- 22
        21204 => X"1E",  -- 30
        21205 => X"31",  -- 49
        21206 => X"4D",  -- 77
        21207 => X"62",  -- 98
        21208 => X"72",  -- 114
        21209 => X"94",  -- 148
        21210 => X"87",  -- 135
        21211 => X"8B",  -- 139
        21212 => X"6F",  -- 111
        21213 => X"5B",  -- 91
        21214 => X"55",  -- 85
        21215 => X"23",  -- 35
        21216 => X"20",  -- 32
        21217 => X"51",  -- 81
        21218 => X"72",  -- 114
        21219 => X"78",  -- 120
        21220 => X"70",  -- 112
        21221 => X"7E",  -- 126
        21222 => X"7F",  -- 127
        21223 => X"7D",  -- 125
        21224 => X"8B",  -- 139
        21225 => X"85",  -- 133
        21226 => X"89",  -- 137
        21227 => X"8B",  -- 139
        21228 => X"99",  -- 153
        21229 => X"91",  -- 145
        21230 => X"8C",  -- 140
        21231 => X"7F",  -- 127
        21232 => X"58",  -- 88
        21233 => X"2A",  -- 42
        21234 => X"07",  -- 7
        21235 => X"06",  -- 6
        21236 => X"10",  -- 16
        21237 => X"0E",  -- 14
        21238 => X"0A",  -- 10
        21239 => X"0C",  -- 12
        21240 => X"09",  -- 9
        21241 => X"1E",  -- 30
        21242 => X"44",  -- 68
        21243 => X"6D",  -- 109
        21244 => X"84",  -- 132
        21245 => X"7E",  -- 126
        21246 => X"6B",  -- 107
        21247 => X"5C",  -- 92
        21248 => X"34",  -- 52
        21249 => X"2F",  -- 47
        21250 => X"20",  -- 32
        21251 => X"13",  -- 19
        21252 => X"20",  -- 32
        21253 => X"45",  -- 69
        21254 => X"66",  -- 102
        21255 => X"74",  -- 116
        21256 => X"64",  -- 100
        21257 => X"3A",  -- 58
        21258 => X"3A",  -- 58
        21259 => X"3A",  -- 58
        21260 => X"4F",  -- 79
        21261 => X"55",  -- 85
        21262 => X"33",  -- 51
        21263 => X"42",  -- 66
        21264 => X"70",  -- 112
        21265 => X"7C",  -- 124
        21266 => X"6F",  -- 111
        21267 => X"5F",  -- 95
        21268 => X"4C",  -- 76
        21269 => X"44",  -- 68
        21270 => X"4D",  -- 77
        21271 => X"46",  -- 70
        21272 => X"66",  -- 102
        21273 => X"6D",  -- 109
        21274 => X"70",  -- 112
        21275 => X"5C",  -- 92
        21276 => X"55",  -- 85
        21277 => X"5E",  -- 94
        21278 => X"56",  -- 86
        21279 => X"5E",  -- 94
        21280 => X"5C",  -- 92
        21281 => X"4C",  -- 76
        21282 => X"43",  -- 67
        21283 => X"32",  -- 50
        21284 => X"3A",  -- 58
        21285 => X"39",  -- 57
        21286 => X"1B",  -- 27
        21287 => X"1F",  -- 31
        21288 => X"67",  -- 103
        21289 => X"B5",  -- 181
        21290 => X"D4",  -- 212
        21291 => X"BE",  -- 190
        21292 => X"C0",  -- 192
        21293 => X"CE",  -- 206
        21294 => X"C8",  -- 200
        21295 => X"C3",  -- 195
        21296 => X"AE",  -- 174
        21297 => X"A3",  -- 163
        21298 => X"98",  -- 152
        21299 => X"96",  -- 150
        21300 => X"94",  -- 148
        21301 => X"8F",  -- 143
        21302 => X"82",  -- 130
        21303 => X"79",  -- 121
        21304 => X"70",  -- 112
        21305 => X"6F",  -- 111
        21306 => X"71",  -- 113
        21307 => X"79",  -- 121
        21308 => X"80",  -- 128
        21309 => X"85",  -- 133
        21310 => X"84",  -- 132
        21311 => X"83",  -- 131
        21312 => X"86",  -- 134
        21313 => X"83",  -- 131
        21314 => X"84",  -- 132
        21315 => X"8B",  -- 139
        21316 => X"97",  -- 151
        21317 => X"A1",  -- 161
        21318 => X"A7",  -- 167
        21319 => X"A9",  -- 169
        21320 => X"9D",  -- 157
        21321 => X"A3",  -- 163
        21322 => X"A9",  -- 169
        21323 => X"A9",  -- 169
        21324 => X"A0",  -- 160
        21325 => X"9E",  -- 158
        21326 => X"A7",  -- 167
        21327 => X"B4",  -- 180
        21328 => X"BA",  -- 186
        21329 => X"BD",  -- 189
        21330 => X"C3",  -- 195
        21331 => X"C6",  -- 198
        21332 => X"C7",  -- 199
        21333 => X"C7",  -- 199
        21334 => X"C6",  -- 198
        21335 => X"C6",  -- 198
        21336 => X"C9",  -- 201
        21337 => X"C7",  -- 199
        21338 => X"C4",  -- 196
        21339 => X"C0",  -- 192
        21340 => X"B3",  -- 179
        21341 => X"9F",  -- 159
        21342 => X"89",  -- 137
        21343 => X"7C",  -- 124
        21344 => X"8B",  -- 139
        21345 => X"A0",  -- 160
        21346 => X"B4",  -- 180
        21347 => X"B9",  -- 185
        21348 => X"B0",  -- 176
        21349 => X"A8",  -- 168
        21350 => X"A5",  -- 165
        21351 => X"A4",  -- 164
        21352 => X"A1",  -- 161
        21353 => X"A1",  -- 161
        21354 => X"A2",  -- 162
        21355 => X"A6",  -- 166
        21356 => X"AA",  -- 170
        21357 => X"AA",  -- 170
        21358 => X"A7",  -- 167
        21359 => X"A4",  -- 164
        21360 => X"9E",  -- 158
        21361 => X"91",  -- 145
        21362 => X"8D",  -- 141
        21363 => X"8C",  -- 140
        21364 => X"8B",  -- 139
        21365 => X"84",  -- 132
        21366 => X"6E",  -- 110
        21367 => X"4F",  -- 79
        21368 => X"3C",  -- 60
        21369 => X"44",  -- 68
        21370 => X"55",  -- 85
        21371 => X"6C",  -- 108
        21372 => X"80",  -- 128
        21373 => X"8C",  -- 140
        21374 => X"92",  -- 146
        21375 => X"96",  -- 150
        21376 => X"93",  -- 147
        21377 => X"8F",  -- 143
        21378 => X"8E",  -- 142
        21379 => X"91",  -- 145
        21380 => X"95",  -- 149
        21381 => X"9C",  -- 156
        21382 => X"9E",  -- 158
        21383 => X"9E",  -- 158
        21384 => X"A1",  -- 161
        21385 => X"A0",  -- 160
        21386 => X"A1",  -- 161
        21387 => X"A5",  -- 165
        21388 => X"AB",  -- 171
        21389 => X"AF",  -- 175
        21390 => X"B2",  -- 178
        21391 => X"B1",  -- 177
        21392 => X"A8",  -- 168
        21393 => X"AE",  -- 174
        21394 => X"A3",  -- 163
        21395 => X"7B",  -- 123
        21396 => X"4B",  -- 75
        21397 => X"2C",  -- 44
        21398 => X"26",  -- 38
        21399 => X"2A",  -- 42
        21400 => X"3A",  -- 58
        21401 => X"58",  -- 88
        21402 => X"78",  -- 120
        21403 => X"86",  -- 134
        21404 => X"8B",  -- 139
        21405 => X"8D",  -- 141
        21406 => X"8D",  -- 141
        21407 => X"8A",  -- 138
        21408 => X"8E",  -- 142
        21409 => X"90",  -- 144
        21410 => X"8E",  -- 142
        21411 => X"89",  -- 137
        21412 => X"85",  -- 133
        21413 => X"88",  -- 136
        21414 => X"92",  -- 146
        21415 => X"9E",  -- 158
        21416 => X"A3",  -- 163
        21417 => X"A6",  -- 166
        21418 => X"AC",  -- 172
        21419 => X"AE",  -- 174
        21420 => X"A7",  -- 167
        21421 => X"9F",  -- 159
        21422 => X"9F",  -- 159
        21423 => X"A3",  -- 163
        21424 => X"A6",  -- 166
        21425 => X"AA",  -- 170
        21426 => X"AF",  -- 175
        21427 => X"B6",  -- 182
        21428 => X"B4",  -- 180
        21429 => X"A8",  -- 168
        21430 => X"92",  -- 146
        21431 => X"80",  -- 128
        21432 => X"8E",  -- 142
        21433 => X"B3",  -- 179
        21434 => X"C5",  -- 197
        21435 => X"BA",  -- 186
        21436 => X"B3",  -- 179
        21437 => X"B9",  -- 185
        21438 => X"BC",  -- 188
        21439 => X"BF",  -- 191
        21440 => X"A5",  -- 165
        21441 => X"A8",  -- 168
        21442 => X"AB",  -- 171
        21443 => X"AD",  -- 173
        21444 => X"AD",  -- 173
        21445 => X"AC",  -- 172
        21446 => X"A8",  -- 168
        21447 => X"A6",  -- 166
        21448 => X"A5",  -- 165
        21449 => X"A5",  -- 165
        21450 => X"A7",  -- 167
        21451 => X"A7",  -- 167
        21452 => X"A7",  -- 167
        21453 => X"A7",  -- 167
        21454 => X"A6",  -- 166
        21455 => X"A6",  -- 166
        21456 => X"A4",  -- 164
        21457 => X"AB",  -- 171
        21458 => X"AB",  -- 171
        21459 => X"A2",  -- 162
        21460 => X"9C",  -- 156
        21461 => X"A0",  -- 160
        21462 => X"9F",  -- 159
        21463 => X"9C",  -- 156
        21464 => X"71",  -- 113
        21465 => X"47",  -- 71
        21466 => X"20",  -- 32
        21467 => X"15",  -- 21
        21468 => X"20",  -- 32
        21469 => X"30",  -- 48
        21470 => X"32",  -- 50
        21471 => X"28",  -- 40
        21472 => X"28",  -- 40
        21473 => X"30",  -- 48
        21474 => X"3B",  -- 59
        21475 => X"3F",  -- 63
        21476 => X"3C",  -- 60
        21477 => X"3E",  -- 62
        21478 => X"42",  -- 66
        21479 => X"44",  -- 68
        21480 => X"24",  -- 36
        21481 => X"2B",  -- 43
        21482 => X"36",  -- 54
        21483 => X"48",  -- 72
        21484 => X"4C",  -- 76
        21485 => X"35",  -- 53
        21486 => X"27",  -- 39
        21487 => X"31",  -- 49
        21488 => X"49",  -- 73
        21489 => X"46",  -- 70
        21490 => X"41",  -- 65
        21491 => X"40",  -- 64
        21492 => X"41",  -- 65
        21493 => X"4B",  -- 75
        21494 => X"63",  -- 99
        21495 => X"7A",  -- 122
        21496 => X"8C",  -- 140
        21497 => X"8B",  -- 139
        21498 => X"79",  -- 121
        21499 => X"4A",  -- 74
        21500 => X"2F",  -- 47
        21501 => X"0D",  -- 13
        21502 => X"0D",  -- 13
        21503 => X"1C",  -- 28
        21504 => X"30",  -- 48
        21505 => X"42",  -- 66
        21506 => X"5C",  -- 92
        21507 => X"79",  -- 121
        21508 => X"8C",  -- 140
        21509 => X"7F",  -- 127
        21510 => X"4D",  -- 77
        21511 => X"1C",  -- 28
        21512 => X"1D",  -- 29
        21513 => X"0C",  -- 12
        21514 => X"09",  -- 9
        21515 => X"05",  -- 5
        21516 => X"09",  -- 9
        21517 => X"17",  -- 23
        21518 => X"10",  -- 16
        21519 => X"16",  -- 22
        21520 => X"1C",  -- 28
        21521 => X"2F",  -- 47
        21522 => X"43",  -- 67
        21523 => X"4F",  -- 79
        21524 => X"5C",  -- 92
        21525 => X"6E",  -- 110
        21526 => X"7E",  -- 126
        21527 => X"88",  -- 136
        21528 => X"8A",  -- 138
        21529 => X"98",  -- 152
        21530 => X"77",  -- 119
        21531 => X"7F",  -- 127
        21532 => X"6F",  -- 111
        21533 => X"5C",  -- 92
        21534 => X"3E",  -- 62
        21535 => X"17",  -- 23
        21536 => X"13",  -- 19
        21537 => X"3D",  -- 61
        21538 => X"6A",  -- 106
        21539 => X"75",  -- 117
        21540 => X"6D",  -- 109
        21541 => X"83",  -- 131
        21542 => X"8F",  -- 143
        21543 => X"85",  -- 133
        21544 => X"92",  -- 146
        21545 => X"80",  -- 128
        21546 => X"78",  -- 120
        21547 => X"7F",  -- 127
        21548 => X"8E",  -- 142
        21549 => X"92",  -- 146
        21550 => X"97",  -- 151
        21551 => X"9C",  -- 156
        21552 => X"9D",  -- 157
        21553 => X"6E",  -- 110
        21554 => X"39",  -- 57
        21555 => X"1E",  -- 30
        21556 => X"10",  -- 16
        21557 => X"07",  -- 7
        21558 => X"08",  -- 8
        21559 => X"0E",  -- 14
        21560 => X"08",  -- 8
        21561 => X"0E",  -- 14
        21562 => X"24",  -- 36
        21563 => X"44",  -- 68
        21564 => X"63",  -- 99
        21565 => X"7A",  -- 122
        21566 => X"7D",  -- 125
        21567 => X"71",  -- 113
        21568 => X"41",  -- 65
        21569 => X"2F",  -- 47
        21570 => X"21",  -- 33
        21571 => X"24",  -- 36
        21572 => X"34",  -- 52
        21573 => X"47",  -- 71
        21574 => X"50",  -- 80
        21575 => X"53",  -- 83
        21576 => X"83",  -- 131
        21577 => X"69",  -- 105
        21578 => X"53",  -- 83
        21579 => X"3F",  -- 63
        21580 => X"51",  -- 81
        21581 => X"63",  -- 99
        21582 => X"4B",  -- 75
        21583 => X"43",  -- 67
        21584 => X"61",  -- 97
        21585 => X"57",  -- 87
        21586 => X"43",  -- 67
        21587 => X"3D",  -- 61
        21588 => X"2D",  -- 45
        21589 => X"12",  -- 18
        21590 => X"11",  -- 17
        21591 => X"10",  -- 16
        21592 => X"1F",  -- 31
        21593 => X"4C",  -- 76
        21594 => X"61",  -- 97
        21595 => X"51",  -- 81
        21596 => X"4F",  -- 79
        21597 => X"3F",  -- 63
        21598 => X"4B",  -- 75
        21599 => X"54",  -- 84
        21600 => X"5C",  -- 92
        21601 => X"47",  -- 71
        21602 => X"4B",  -- 75
        21603 => X"3F",  -- 63
        21604 => X"3C",  -- 60
        21605 => X"2B",  -- 43
        21606 => X"1D",  -- 29
        21607 => X"5C",  -- 92
        21608 => X"BE",  -- 190
        21609 => X"C4",  -- 196
        21610 => X"BD",  -- 189
        21611 => X"B9",  -- 185
        21612 => X"BF",  -- 191
        21613 => X"BD",  -- 189
        21614 => X"BB",  -- 187
        21615 => X"CB",  -- 203
        21616 => X"BD",  -- 189
        21617 => X"A2",  -- 162
        21618 => X"86",  -- 134
        21619 => X"80",  -- 128
        21620 => X"8A",  -- 138
        21621 => X"90",  -- 144
        21622 => X"8C",  -- 140
        21623 => X"85",  -- 133
        21624 => X"7B",  -- 123
        21625 => X"76",  -- 118
        21626 => X"72",  -- 114
        21627 => X"71",  -- 113
        21628 => X"78",  -- 120
        21629 => X"81",  -- 129
        21630 => X"86",  -- 134
        21631 => X"8A",  -- 138
        21632 => X"86",  -- 134
        21633 => X"83",  -- 131
        21634 => X"82",  -- 130
        21635 => X"88",  -- 136
        21636 => X"94",  -- 148
        21637 => X"A0",  -- 160
        21638 => X"A6",  -- 166
        21639 => X"A9",  -- 169
        21640 => X"A1",  -- 161
        21641 => X"A5",  -- 165
        21642 => X"A9",  -- 169
        21643 => X"A7",  -- 167
        21644 => X"A3",  -- 163
        21645 => X"A1",  -- 161
        21646 => X"AC",  -- 172
        21647 => X"BA",  -- 186
        21648 => X"C0",  -- 192
        21649 => X"BF",  -- 191
        21650 => X"BF",  -- 191
        21651 => X"BE",  -- 190
        21652 => X"BF",  -- 191
        21653 => X"C3",  -- 195
        21654 => X"C8",  -- 200
        21655 => X"CD",  -- 205
        21656 => X"CF",  -- 207
        21657 => X"CC",  -- 204
        21658 => X"C9",  -- 201
        21659 => X"C6",  -- 198
        21660 => X"BD",  -- 189
        21661 => X"A5",  -- 165
        21662 => X"88",  -- 136
        21663 => X"72",  -- 114
        21664 => X"7E",  -- 126
        21665 => X"96",  -- 150
        21666 => X"AE",  -- 174
        21667 => X"B6",  -- 182
        21668 => X"B1",  -- 177
        21669 => X"A8",  -- 168
        21670 => X"A1",  -- 161
        21671 => X"9B",  -- 155
        21672 => X"9B",  -- 155
        21673 => X"9E",  -- 158
        21674 => X"A1",  -- 161
        21675 => X"A6",  -- 166
        21676 => X"AA",  -- 170
        21677 => X"AA",  -- 170
        21678 => X"A7",  -- 167
        21679 => X"A4",  -- 164
        21680 => X"98",  -- 152
        21681 => X"91",  -- 145
        21682 => X"90",  -- 144
        21683 => X"91",  -- 145
        21684 => X"8A",  -- 138
        21685 => X"7D",  -- 125
        21686 => X"63",  -- 99
        21687 => X"46",  -- 70
        21688 => X"43",  -- 67
        21689 => X"4B",  -- 75
        21690 => X"5B",  -- 91
        21691 => X"6E",  -- 110
        21692 => X"7C",  -- 124
        21693 => X"87",  -- 135
        21694 => X"8D",  -- 141
        21695 => X"92",  -- 146
        21696 => X"95",  -- 149
        21697 => X"93",  -- 147
        21698 => X"92",  -- 146
        21699 => X"92",  -- 146
        21700 => X"95",  -- 149
        21701 => X"9A",  -- 154
        21702 => X"A1",  -- 161
        21703 => X"A5",  -- 165
        21704 => X"9E",  -- 158
        21705 => X"A0",  -- 160
        21706 => X"A1",  -- 161
        21707 => X"A3",  -- 163
        21708 => X"A8",  -- 168
        21709 => X"AD",  -- 173
        21710 => X"B1",  -- 177
        21711 => X"B4",  -- 180
        21712 => X"BC",  -- 188
        21713 => X"B3",  -- 179
        21714 => X"AB",  -- 171
        21715 => X"96",  -- 150
        21716 => X"68",  -- 104
        21717 => X"35",  -- 53
        21718 => X"22",  -- 34
        21719 => X"2C",  -- 44
        21720 => X"42",  -- 66
        21721 => X"61",  -- 97
        21722 => X"81",  -- 129
        21723 => X"8F",  -- 143
        21724 => X"91",  -- 145
        21725 => X"8F",  -- 143
        21726 => X"8D",  -- 141
        21727 => X"88",  -- 136
        21728 => X"90",  -- 144
        21729 => X"81",  -- 129
        21730 => X"70",  -- 112
        21731 => X"6C",  -- 108
        21732 => X"72",  -- 114
        21733 => X"80",  -- 128
        21734 => X"90",  -- 144
        21735 => X"9C",  -- 156
        21736 => X"A6",  -- 166
        21737 => X"A8",  -- 168
        21738 => X"AE",  -- 174
        21739 => X"AF",  -- 175
        21740 => X"AB",  -- 171
        21741 => X"A2",  -- 162
        21742 => X"9D",  -- 157
        21743 => X"9E",  -- 158
        21744 => X"9E",  -- 158
        21745 => X"A5",  -- 165
        21746 => X"AC",  -- 172
        21747 => X"AF",  -- 175
        21748 => X"B0",  -- 176
        21749 => X"A6",  -- 166
        21750 => X"90",  -- 144
        21751 => X"7B",  -- 123
        21752 => X"89",  -- 137
        21753 => X"B6",  -- 182
        21754 => X"CB",  -- 203
        21755 => X"BB",  -- 187
        21756 => X"B0",  -- 176
        21757 => X"B2",  -- 178
        21758 => X"B5",  -- 181
        21759 => X"B6",  -- 182
        21760 => X"AC",  -- 172
        21761 => X"AB",  -- 171
        21762 => X"AC",  -- 172
        21763 => X"AB",  -- 171
        21764 => X"AB",  -- 171
        21765 => X"AA",  -- 170
        21766 => X"AB",  -- 171
        21767 => X"AA",  -- 170
        21768 => X"A8",  -- 168
        21769 => X"A8",  -- 168
        21770 => X"A7",  -- 167
        21771 => X"A7",  -- 167
        21772 => X"A8",  -- 168
        21773 => X"A8",  -- 168
        21774 => X"A8",  -- 168
        21775 => X"A8",  -- 168
        21776 => X"AC",  -- 172
        21777 => X"A7",  -- 167
        21778 => X"A6",  -- 166
        21779 => X"AB",  -- 171
        21780 => X"AC",  -- 172
        21781 => X"A6",  -- 166
        21782 => X"9E",  -- 158
        21783 => X"9B",  -- 155
        21784 => X"AA",  -- 170
        21785 => X"83",  -- 131
        21786 => X"57",  -- 87
        21787 => X"33",  -- 51
        21788 => X"1B",  -- 27
        21789 => X"1B",  -- 27
        21790 => X"29",  -- 41
        21791 => X"34",  -- 52
        21792 => X"2A",  -- 42
        21793 => X"36",  -- 54
        21794 => X"39",  -- 57
        21795 => X"35",  -- 53
        21796 => X"39",  -- 57
        21797 => X"3B",  -- 59
        21798 => X"2E",  -- 46
        21799 => X"1F",  -- 31
        21800 => X"18",  -- 24
        21801 => X"1C",  -- 28
        21802 => X"1A",  -- 26
        21803 => X"1F",  -- 31
        21804 => X"25",  -- 37
        21805 => X"23",  -- 35
        21806 => X"2A",  -- 42
        21807 => X"3A",  -- 58
        21808 => X"3D",  -- 61
        21809 => X"25",  -- 37
        21810 => X"2D",  -- 45
        21811 => X"51",  -- 81
        21812 => X"59",  -- 89
        21813 => X"4D",  -- 77
        21814 => X"68",  -- 104
        21815 => X"9B",  -- 155
        21816 => X"91",  -- 145
        21817 => X"7B",  -- 123
        21818 => X"64",  -- 100
        21819 => X"31",  -- 49
        21820 => X"17",  -- 23
        21821 => X"14",  -- 20
        21822 => X"2B",  -- 43
        21823 => X"29",  -- 41
        21824 => X"22",  -- 34
        21825 => X"42",  -- 66
        21826 => X"72",  -- 114
        21827 => X"8E",  -- 142
        21828 => X"85",  -- 133
        21829 => X"5B",  -- 91
        21830 => X"29",  -- 41
        21831 => X"0B",  -- 11
        21832 => X"07",  -- 7
        21833 => X"0A",  -- 10
        21834 => X"04",  -- 4
        21835 => X"04",  -- 4
        21836 => X"09",  -- 9
        21837 => X"11",  -- 17
        21838 => X"30",  -- 48
        21839 => X"38",  -- 56
        21840 => X"51",  -- 81
        21841 => X"64",  -- 100
        21842 => X"7B",  -- 123
        21843 => X"8A",  -- 138
        21844 => X"92",  -- 146
        21845 => X"96",  -- 150
        21846 => X"95",  -- 149
        21847 => X"94",  -- 148
        21848 => X"9B",  -- 155
        21849 => X"93",  -- 147
        21850 => X"7F",  -- 127
        21851 => X"83",  -- 131
        21852 => X"71",  -- 113
        21853 => X"54",  -- 84
        21854 => X"1C",  -- 28
        21855 => X"0C",  -- 12
        21856 => X"0B",  -- 11
        21857 => X"21",  -- 33
        21858 => X"56",  -- 86
        21859 => X"72",  -- 114
        21860 => X"74",  -- 116
        21861 => X"7C",  -- 124
        21862 => X"8D",  -- 141
        21863 => X"89",  -- 137
        21864 => X"82",  -- 130
        21865 => X"75",  -- 117
        21866 => X"6F",  -- 111
        21867 => X"80",  -- 128
        21868 => X"8A",  -- 138
        21869 => X"8E",  -- 142
        21870 => X"8F",  -- 143
        21871 => X"9A",  -- 154
        21872 => X"A0",  -- 160
        21873 => X"97",  -- 151
        21874 => X"7B",  -- 123
        21875 => X"49",  -- 73
        21876 => X"1C",  -- 28
        21877 => X"08",  -- 8
        21878 => X"07",  -- 7
        21879 => X"0D",  -- 13
        21880 => X"04",  -- 4
        21881 => X"07",  -- 7
        21882 => X"16",  -- 22
        21883 => X"26",  -- 38
        21884 => X"40",  -- 64
        21885 => X"68",  -- 104
        21886 => X"81",  -- 129
        21887 => X"7A",  -- 122
        21888 => X"6C",  -- 108
        21889 => X"4A",  -- 74
        21890 => X"3A",  -- 58
        21891 => X"44",  -- 68
        21892 => X"4A",  -- 74
        21893 => X"42",  -- 66
        21894 => X"44",  -- 68
        21895 => X"52",  -- 82
        21896 => X"6F",  -- 111
        21897 => X"92",  -- 146
        21898 => X"89",  -- 137
        21899 => X"70",  -- 112
        21900 => X"55",  -- 85
        21901 => X"4A",  -- 74
        21902 => X"67",  -- 103
        21903 => X"77",  -- 119
        21904 => X"43",  -- 67
        21905 => X"46",  -- 70
        21906 => X"3F",  -- 63
        21907 => X"3A",  -- 58
        21908 => X"24",  -- 36
        21909 => X"0E",  -- 14
        21910 => X"1C",  -- 28
        21911 => X"2B",  -- 43
        21912 => X"17",  -- 23
        21913 => X"2F",  -- 47
        21914 => X"32",  -- 50
        21915 => X"21",  -- 33
        21916 => X"29",  -- 41
        21917 => X"1A",  -- 26
        21918 => X"3C",  -- 60
        21919 => X"4F",  -- 79
        21920 => X"56",  -- 86
        21921 => X"4F",  -- 79
        21922 => X"5D",  -- 93
        21923 => X"47",  -- 71
        21924 => X"2E",  -- 46
        21925 => X"1D",  -- 29
        21926 => X"34",  -- 52
        21927 => X"9C",  -- 156
        21928 => X"BE",  -- 190
        21929 => X"B3",  -- 179
        21930 => X"B2",  -- 178
        21931 => X"AC",  -- 172
        21932 => X"A4",  -- 164
        21933 => X"AD",  -- 173
        21934 => X"BA",  -- 186
        21935 => X"B8",  -- 184
        21936 => X"B4",  -- 180
        21937 => X"A0",  -- 160
        21938 => X"88",  -- 136
        21939 => X"79",  -- 121
        21940 => X"6F",  -- 111
        21941 => X"6F",  -- 111
        21942 => X"77",  -- 119
        21943 => X"81",  -- 129
        21944 => X"74",  -- 116
        21945 => X"72",  -- 114
        21946 => X"71",  -- 113
        21947 => X"76",  -- 118
        21948 => X"7C",  -- 124
        21949 => X"83",  -- 131
        21950 => X"88",  -- 136
        21951 => X"8A",  -- 138
        21952 => X"87",  -- 135
        21953 => X"88",  -- 136
        21954 => X"89",  -- 137
        21955 => X"8C",  -- 140
        21956 => X"92",  -- 146
        21957 => X"98",  -- 152
        21958 => X"A2",  -- 162
        21959 => X"A7",  -- 167
        21960 => X"A3",  -- 163
        21961 => X"A0",  -- 160
        21962 => X"9F",  -- 159
        21963 => X"A1",  -- 161
        21964 => X"A4",  -- 164
        21965 => X"A9",  -- 169
        21966 => X"B6",  -- 182
        21967 => X"C0",  -- 192
        21968 => X"C0",  -- 192
        21969 => X"BF",  -- 191
        21970 => X"BD",  -- 189
        21971 => X"BB",  -- 187
        21972 => X"BB",  -- 187
        21973 => X"C0",  -- 192
        21974 => X"C9",  -- 201
        21975 => X"CE",  -- 206
        21976 => X"CF",  -- 207
        21977 => X"CD",  -- 205
        21978 => X"CC",  -- 204
        21979 => X"C8",  -- 200
        21980 => X"BD",  -- 189
        21981 => X"A9",  -- 169
        21982 => X"8A",  -- 138
        21983 => X"74",  -- 116
        21984 => X"81",  -- 129
        21985 => X"91",  -- 145
        21986 => X"A3",  -- 163
        21987 => X"AD",  -- 173
        21988 => X"B1",  -- 177
        21989 => X"AF",  -- 175
        21990 => X"A8",  -- 168
        21991 => X"9F",  -- 159
        21992 => X"9E",  -- 158
        21993 => X"A0",  -- 160
        21994 => X"A3",  -- 163
        21995 => X"A7",  -- 167
        21996 => X"A7",  -- 167
        21997 => X"A4",  -- 164
        21998 => X"A0",  -- 160
        21999 => X"9C",  -- 156
        22000 => X"91",  -- 145
        22001 => X"8E",  -- 142
        22002 => X"92",  -- 146
        22003 => X"90",  -- 144
        22004 => X"85",  -- 133
        22005 => X"79",  -- 121
        22006 => X"63",  -- 99
        22007 => X"4B",  -- 75
        22008 => X"4A",  -- 74
        22009 => X"4A",  -- 74
        22010 => X"52",  -- 82
        22011 => X"65",  -- 101
        22012 => X"80",  -- 128
        22013 => X"8F",  -- 143
        22014 => X"8E",  -- 142
        22015 => X"87",  -- 135
        22016 => X"8F",  -- 143
        22017 => X"97",  -- 151
        22018 => X"A0",  -- 160
        22019 => X"A4",  -- 164
        22020 => X"A1",  -- 161
        22021 => X"A0",  -- 160
        22022 => X"A1",  -- 161
        22023 => X"A3",  -- 163
        22024 => X"A2",  -- 162
        22025 => X"A3",  -- 163
        22026 => X"A5",  -- 165
        22027 => X"A9",  -- 169
        22028 => X"AC",  -- 172
        22029 => X"B2",  -- 178
        22030 => X"B6",  -- 182
        22031 => X"BA",  -- 186
        22032 => X"BC",  -- 188
        22033 => X"B5",  -- 181
        22034 => X"AC",  -- 172
        22035 => X"8F",  -- 143
        22036 => X"54",  -- 84
        22037 => X"1F",  -- 31
        22038 => X"1D",  -- 29
        22039 => X"37",  -- 55
        22040 => X"5C",  -- 92
        22041 => X"72",  -- 114
        22042 => X"86",  -- 134
        22043 => X"8C",  -- 140
        22044 => X"8C",  -- 140
        22045 => X"90",  -- 144
        22046 => X"94",  -- 148
        22047 => X"94",  -- 148
        22048 => X"88",  -- 136
        22049 => X"72",  -- 114
        22050 => X"63",  -- 99
        22051 => X"67",  -- 103
        22052 => X"79",  -- 121
        22053 => X"8B",  -- 139
        22054 => X"9A",  -- 154
        22055 => X"A2",  -- 162
        22056 => X"AE",  -- 174
        22057 => X"AD",  -- 173
        22058 => X"B0",  -- 176
        22059 => X"B6",  -- 182
        22060 => X"B5",  -- 181
        22061 => X"A9",  -- 169
        22062 => X"9C",  -- 156
        22063 => X"96",  -- 150
        22064 => X"99",  -- 153
        22065 => X"A1",  -- 161
        22066 => X"AA",  -- 170
        22067 => X"AC",  -- 172
        22068 => X"AD",  -- 173
        22069 => X"A6",  -- 166
        22070 => X"8F",  -- 143
        22071 => X"75",  -- 117
        22072 => X"8B",  -- 139
        22073 => X"B7",  -- 183
        22074 => X"C8",  -- 200
        22075 => X"B6",  -- 182
        22076 => X"A5",  -- 165
        22077 => X"A6",  -- 166
        22078 => X"AA",  -- 170
        22079 => X"AB",  -- 171
        22080 => X"B4",  -- 180
        22081 => X"B3",  -- 179
        22082 => X"B2",  -- 178
        22083 => X"B1",  -- 177
        22084 => X"AF",  -- 175
        22085 => X"AE",  -- 174
        22086 => X"AF",  -- 175
        22087 => X"B0",  -- 176
        22088 => X"AE",  -- 174
        22089 => X"AC",  -- 172
        22090 => X"A8",  -- 168
        22091 => X"A7",  -- 167
        22092 => X"A9",  -- 169
        22093 => X"A9",  -- 169
        22094 => X"A9",  -- 169
        22095 => X"A9",  -- 169
        22096 => X"AA",  -- 170
        22097 => X"A9",  -- 169
        22098 => X"A5",  -- 165
        22099 => X"A5",  -- 165
        22100 => X"A8",  -- 168
        22101 => X"AB",  -- 171
        22102 => X"A4",  -- 164
        22103 => X"9A",  -- 154
        22104 => X"9C",  -- 156
        22105 => X"9D",  -- 157
        22106 => X"95",  -- 149
        22107 => X"76",  -- 118
        22108 => X"48",  -- 72
        22109 => X"26",  -- 38
        22110 => X"21",  -- 33
        22111 => X"2F",  -- 47
        22112 => X"3A",  -- 58
        22113 => X"50",  -- 80
        22114 => X"54",  -- 84
        22115 => X"4E",  -- 78
        22116 => X"54",  -- 84
        22117 => X"55",  -- 85
        22118 => X"3F",  -- 63
        22119 => X"2C",  -- 44
        22120 => X"4B",  -- 75
        22121 => X"51",  -- 81
        22122 => X"4F",  -- 79
        22123 => X"4E",  -- 78
        22124 => X"51",  -- 81
        22125 => X"48",  -- 72
        22126 => X"39",  -- 57
        22127 => X"34",  -- 52
        22128 => X"2B",  -- 43
        22129 => X"30",  -- 48
        22130 => X"3C",  -- 60
        22131 => X"4C",  -- 76
        22132 => X"58",  -- 88
        22133 => X"66",  -- 102
        22134 => X"7B",  -- 123
        22135 => X"8E",  -- 142
        22136 => X"79",  -- 121
        22137 => X"58",  -- 88
        22138 => X"46",  -- 70
        22139 => X"23",  -- 35
        22140 => X"1B",  -- 27
        22141 => X"2B",  -- 43
        22142 => X"48",  -- 72
        22143 => X"37",  -- 55
        22144 => X"41",  -- 65
        22145 => X"58",  -- 88
        22146 => X"77",  -- 119
        22147 => X"7E",  -- 126
        22148 => X"5C",  -- 92
        22149 => X"2B",  -- 43
        22150 => X"0E",  -- 14
        22151 => X"08",  -- 8
        22152 => X"09",  -- 9
        22153 => X"1C",  -- 28
        22154 => X"1E",  -- 30
        22155 => X"29",  -- 41
        22156 => X"38",  -- 56
        22157 => X"41",  -- 65
        22158 => X"73",  -- 115
        22159 => X"7C",  -- 124
        22160 => X"8A",  -- 138
        22161 => X"92",  -- 146
        22162 => X"9D",  -- 157
        22163 => X"A2",  -- 162
        22164 => X"9D",  -- 157
        22165 => X"96",  -- 150
        22166 => X"96",  -- 150
        22167 => X"9C",  -- 156
        22168 => X"99",  -- 153
        22169 => X"8F",  -- 143
        22170 => X"90",  -- 144
        22171 => X"8B",  -- 139
        22172 => X"69",  -- 105
        22173 => X"38",  -- 56
        22174 => X"0B",  -- 11
        22175 => X"0E",  -- 14
        22176 => X"25",  -- 37
        22177 => X"0A",  -- 10
        22178 => X"26",  -- 38
        22179 => X"60",  -- 96
        22180 => X"88",  -- 136
        22181 => X"87",  -- 135
        22182 => X"84",  -- 132
        22183 => X"76",  -- 118
        22184 => X"59",  -- 89
        22185 => X"4E",  -- 78
        22186 => X"47",  -- 71
        22187 => X"57",  -- 87
        22188 => X"5C",  -- 92
        22189 => X"63",  -- 99
        22190 => X"66",  -- 102
        22191 => X"75",  -- 117
        22192 => X"8B",  -- 139
        22193 => X"98",  -- 152
        22194 => X"92",  -- 146
        22195 => X"6F",  -- 111
        22196 => X"4E",  -- 78
        22197 => X"3B",  -- 59
        22198 => X"20",  -- 32
        22199 => X"06",  -- 6
        22200 => X"03",  -- 3
        22201 => X"03",  -- 3
        22202 => X"0A",  -- 10
        22203 => X"10",  -- 16
        22204 => X"1C",  -- 28
        22205 => X"48",  -- 72
        22206 => X"74",  -- 116
        22207 => X"7C",  -- 124
        22208 => X"7C",  -- 124
        22209 => X"7B",  -- 123
        22210 => X"68",  -- 104
        22211 => X"48",  -- 72
        22212 => X"34",  -- 52
        22213 => X"37",  -- 55
        22214 => X"44",  -- 68
        22215 => X"4B",  -- 75
        22216 => X"57",  -- 87
        22217 => X"81",  -- 129
        22218 => X"83",  -- 131
        22219 => X"94",  -- 148
        22220 => X"7D",  -- 125
        22221 => X"54",  -- 84
        22222 => X"67",  -- 103
        22223 => X"6F",  -- 111
        22224 => X"6F",  -- 111
        22225 => X"5F",  -- 95
        22226 => X"3D",  -- 61
        22227 => X"36",  -- 54
        22228 => X"40",  -- 64
        22229 => X"43",  -- 67
        22230 => X"36",  -- 54
        22231 => X"15",  -- 21
        22232 => X"1E",  -- 30
        22233 => X"16",  -- 22
        22234 => X"0E",  -- 14
        22235 => X"0A",  -- 10
        22236 => X"21",  -- 33
        22237 => X"1F",  -- 31
        22238 => X"32",  -- 50
        22239 => X"38",  -- 56
        22240 => X"51",  -- 81
        22241 => X"62",  -- 98
        22242 => X"74",  -- 116
        22243 => X"4D",  -- 77
        22244 => X"1B",  -- 27
        22245 => X"10",  -- 16
        22246 => X"40",  -- 64
        22247 => X"A5",  -- 165
        22248 => X"BC",  -- 188
        22249 => X"AE",  -- 174
        22250 => X"AB",  -- 171
        22251 => X"9B",  -- 155
        22252 => X"8B",  -- 139
        22253 => X"A2",  -- 162
        22254 => X"B4",  -- 180
        22255 => X"A4",  -- 164
        22256 => X"9C",  -- 156
        22257 => X"8E",  -- 142
        22258 => X"7E",  -- 126
        22259 => X"6E",  -- 110
        22260 => X"5D",  -- 93
        22261 => X"4E",  -- 78
        22262 => X"4C",  -- 76
        22263 => X"51",  -- 81
        22264 => X"4C",  -- 76
        22265 => X"54",  -- 84
        22266 => X"5F",  -- 95
        22267 => X"6D",  -- 109
        22268 => X"79",  -- 121
        22269 => X"80",  -- 128
        22270 => X"80",  -- 128
        22271 => X"7F",  -- 127
        22272 => X"8D",  -- 141
        22273 => X"90",  -- 144
        22274 => X"94",  -- 148
        22275 => X"95",  -- 149
        22276 => X"94",  -- 148
        22277 => X"9A",  -- 154
        22278 => X"A3",  -- 163
        22279 => X"AD",  -- 173
        22280 => X"B1",  -- 177
        22281 => X"A8",  -- 168
        22282 => X"A2",  -- 162
        22283 => X"A5",  -- 165
        22284 => X"AA",  -- 170
        22285 => X"AF",  -- 175
        22286 => X"B7",  -- 183
        22287 => X"BC",  -- 188
        22288 => X"C2",  -- 194
        22289 => X"C2",  -- 194
        22290 => X"C4",  -- 196
        22291 => X"C5",  -- 197
        22292 => X"C6",  -- 198
        22293 => X"C8",  -- 200
        22294 => X"CB",  -- 203
        22295 => X"CE",  -- 206
        22296 => X"CB",  -- 203
        22297 => X"CC",  -- 204
        22298 => X"CA",  -- 202
        22299 => X"C6",  -- 198
        22300 => X"BC",  -- 188
        22301 => X"AD",  -- 173
        22302 => X"96",  -- 150
        22303 => X"83",  -- 131
        22304 => X"88",  -- 136
        22305 => X"8C",  -- 140
        22306 => X"94",  -- 148
        22307 => X"9D",  -- 157
        22308 => X"A9",  -- 169
        22309 => X"AF",  -- 175
        22310 => X"AD",  -- 173
        22311 => X"A7",  -- 167
        22312 => X"A7",  -- 167
        22313 => X"A7",  -- 167
        22314 => X"A7",  -- 167
        22315 => X"A6",  -- 166
        22316 => X"A4",  -- 164
        22317 => X"A0",  -- 160
        22318 => X"9B",  -- 155
        22319 => X"97",  -- 151
        22320 => X"96",  -- 150
        22321 => X"90",  -- 144
        22322 => X"93",  -- 147
        22323 => X"90",  -- 144
        22324 => X"89",  -- 137
        22325 => X"81",  -- 129
        22326 => X"74",  -- 116
        22327 => X"60",  -- 96
        22328 => X"3E",  -- 62
        22329 => X"44",  -- 68
        22330 => X"4E",  -- 78
        22331 => X"61",  -- 97
        22332 => X"78",  -- 120
        22333 => X"8C",  -- 140
        22334 => X"92",  -- 146
        22335 => X"92",  -- 146
        22336 => X"93",  -- 147
        22337 => X"98",  -- 152
        22338 => X"9F",  -- 159
        22339 => X"9F",  -- 159
        22340 => X"9D",  -- 157
        22341 => X"9D",  -- 157
        22342 => X"A2",  -- 162
        22343 => X"A6",  -- 166
        22344 => X"A6",  -- 166
        22345 => X"A6",  -- 166
        22346 => X"A9",  -- 169
        22347 => X"AC",  -- 172
        22348 => X"B2",  -- 178
        22349 => X"B6",  -- 182
        22350 => X"B9",  -- 185
        22351 => X"BA",  -- 186
        22352 => X"B7",  -- 183
        22353 => X"B6",  -- 182
        22354 => X"A8",  -- 168
        22355 => X"81",  -- 129
        22356 => X"46",  -- 70
        22357 => X"21",  -- 33
        22358 => X"23",  -- 35
        22359 => X"36",  -- 54
        22360 => X"65",  -- 101
        22361 => X"78",  -- 120
        22362 => X"88",  -- 136
        22363 => X"8B",  -- 139
        22364 => X"8B",  -- 139
        22365 => X"8E",  -- 142
        22366 => X"90",  -- 144
        22367 => X"8E",  -- 142
        22368 => X"87",  -- 135
        22369 => X"7B",  -- 123
        22370 => X"76",  -- 118
        22371 => X"84",  -- 132
        22372 => X"96",  -- 150
        22373 => X"A1",  -- 161
        22374 => X"A3",  -- 163
        22375 => X"A3",  -- 163
        22376 => X"AE",  -- 174
        22377 => X"AB",  -- 171
        22378 => X"AF",  -- 175
        22379 => X"B6",  -- 182
        22380 => X"B6",  -- 182
        22381 => X"AA",  -- 170
        22382 => X"99",  -- 153
        22383 => X"90",  -- 144
        22384 => X"9E",  -- 158
        22385 => X"A7",  -- 167
        22386 => X"AC",  -- 172
        22387 => X"AD",  -- 173
        22388 => X"B0",  -- 176
        22389 => X"AC",  -- 172
        22390 => X"8F",  -- 143
        22391 => X"71",  -- 113
        22392 => X"83",  -- 131
        22393 => X"AA",  -- 170
        22394 => X"BA",  -- 186
        22395 => X"AA",  -- 170
        22396 => X"9C",  -- 156
        22397 => X"A0",  -- 160
        22398 => X"A9",  -- 169
        22399 => X"B2",  -- 178
        22400 => X"B4",  -- 180
        22401 => X"B4",  -- 180
        22402 => X"B4",  -- 180
        22403 => X"B3",  -- 179
        22404 => X"B2",  -- 178
        22405 => X"B0",  -- 176
        22406 => X"AF",  -- 175
        22407 => X"AE",  -- 174
        22408 => X"AC",  -- 172
        22409 => X"A8",  -- 168
        22410 => X"A3",  -- 163
        22411 => X"A1",  -- 161
        22412 => X"A2",  -- 162
        22413 => X"A3",  -- 163
        22414 => X"A3",  -- 163
        22415 => X"A3",  -- 163
        22416 => X"9E",  -- 158
        22417 => X"9F",  -- 159
        22418 => X"9A",  -- 154
        22419 => X"93",  -- 147
        22420 => X"8F",  -- 143
        22421 => X"96",  -- 150
        22422 => X"9D",  -- 157
        22423 => X"A0",  -- 160
        22424 => X"A0",  -- 160
        22425 => X"9B",  -- 155
        22426 => X"8A",  -- 138
        22427 => X"83",  -- 131
        22428 => X"79",  -- 121
        22429 => X"4B",  -- 75
        22430 => X"16",  -- 22
        22431 => X"02",  -- 2
        22432 => X"38",  -- 56
        22433 => X"45",  -- 69
        22434 => X"3F",  -- 63
        22435 => X"36",  -- 54
        22436 => X"45",  -- 69
        22437 => X"57",  -- 87
        22438 => X"66",  -- 102
        22439 => X"75",  -- 117
        22440 => X"6B",  -- 107
        22441 => X"67",  -- 103
        22442 => X"57",  -- 87
        22443 => X"4A",  -- 74
        22444 => X"46",  -- 70
        22445 => X"3E",  -- 62
        22446 => X"3B",  -- 59
        22447 => X"42",  -- 66
        22448 => X"36",  -- 54
        22449 => X"4A",  -- 74
        22450 => X"4A",  -- 74
        22451 => X"3D",  -- 61
        22452 => X"56",  -- 86
        22453 => X"81",  -- 129
        22454 => X"82",  -- 130
        22455 => X"5E",  -- 94
        22456 => X"4F",  -- 79
        22457 => X"36",  -- 54
        22458 => X"26",  -- 38
        22459 => X"1C",  -- 28
        22460 => X"33",  -- 51
        22461 => X"49",  -- 73
        22462 => X"5C",  -- 92
        22463 => X"52",  -- 82
        22464 => X"6F",  -- 111
        22465 => X"6D",  -- 109
        22466 => X"67",  -- 103
        22467 => X"5B",  -- 91
        22468 => X"3E",  -- 62
        22469 => X"21",  -- 33
        22470 => X"16",  -- 22
        22471 => X"18",  -- 24
        22472 => X"3D",  -- 61
        22473 => X"4C",  -- 76
        22474 => X"62",  -- 98
        22475 => X"67",  -- 103
        22476 => X"79",  -- 121
        22477 => X"7D",  -- 125
        22478 => X"97",  -- 151
        22479 => X"9B",  -- 155
        22480 => X"94",  -- 148
        22481 => X"92",  -- 146
        22482 => X"91",  -- 145
        22483 => X"8C",  -- 140
        22484 => X"7E",  -- 126
        22485 => X"79",  -- 121
        22486 => X"89",  -- 137
        22487 => X"A3",  -- 163
        22488 => X"90",  -- 144
        22489 => X"8D",  -- 141
        22490 => X"8A",  -- 138
        22491 => X"7A",  -- 122
        22492 => X"4F",  -- 79
        22493 => X"19",  -- 25
        22494 => X"12",  -- 18
        22495 => X"1B",  -- 27
        22496 => X"38",  -- 56
        22497 => X"06",  -- 6
        22498 => X"07",  -- 7
        22499 => X"34",  -- 52
        22500 => X"7D",  -- 125
        22501 => X"8C",  -- 140
        22502 => X"81",  -- 129
        22503 => X"62",  -- 98
        22504 => X"3B",  -- 59
        22505 => X"2C",  -- 44
        22506 => X"18",  -- 24
        22507 => X"20",  -- 32
        22508 => X"1C",  -- 28
        22509 => X"29",  -- 41
        22510 => X"2D",  -- 45
        22511 => X"3B",  -- 59
        22512 => X"78",  -- 120
        22513 => X"86",  -- 134
        22514 => X"8B",  -- 139
        22515 => X"85",  -- 133
        22516 => X"84",  -- 132
        22517 => X"7D",  -- 125
        22518 => X"56",  -- 86
        22519 => X"2A",  -- 42
        22520 => X"1E",  -- 30
        22521 => X"10",  -- 16
        22522 => X"14",  -- 20
        22523 => X"16",  -- 22
        22524 => X"0F",  -- 15
        22525 => X"27",  -- 39
        22526 => X"56",  -- 86
        22527 => X"6D",  -- 109
        22528 => X"7C",  -- 124
        22529 => X"91",  -- 145
        22530 => X"89",  -- 137
        22531 => X"59",  -- 89
        22532 => X"2F",  -- 47
        22533 => X"28",  -- 40
        22534 => X"2D",  -- 45
        22535 => X"2E",  -- 46
        22536 => X"37",  -- 55
        22537 => X"48",  -- 72
        22538 => X"53",  -- 83
        22539 => X"81",  -- 129
        22540 => X"9C",  -- 156
        22541 => X"85",  -- 133
        22542 => X"76",  -- 118
        22543 => X"65",  -- 101
        22544 => X"72",  -- 114
        22545 => X"83",  -- 131
        22546 => X"76",  -- 118
        22547 => X"57",  -- 87
        22548 => X"31",  -- 49
        22549 => X"1D",  -- 29
        22550 => X"27",  -- 39
        22551 => X"29",  -- 41
        22552 => X"0B",  -- 11
        22553 => X"05",  -- 5
        22554 => X"12",  -- 18
        22555 => X"15",  -- 21
        22556 => X"21",  -- 33
        22557 => X"21",  -- 33
        22558 => X"22",  -- 34
        22559 => X"1C",  -- 28
        22560 => X"4C",  -- 76
        22561 => X"67",  -- 103
        22562 => X"7E",  -- 126
        22563 => X"63",  -- 99
        22564 => X"29",  -- 41
        22565 => X"14",  -- 20
        22566 => X"4C",  -- 76
        22567 => X"9D",  -- 157
        22568 => X"C0",  -- 192
        22569 => X"AE",  -- 174
        22570 => X"9B",  -- 155
        22571 => X"8C",  -- 140
        22572 => X"86",  -- 134
        22573 => X"91",  -- 145
        22574 => X"9E",  -- 158
        22575 => X"A1",  -- 161
        22576 => X"9A",  -- 154
        22577 => X"80",  -- 128
        22578 => X"69",  -- 105
        22579 => X"65",  -- 101
        22580 => X"61",  -- 97
        22581 => X"52",  -- 82
        22582 => X"3E",  -- 62
        22583 => X"32",  -- 50
        22584 => X"32",  -- 50
        22585 => X"38",  -- 56
        22586 => X"45",  -- 69
        22587 => X"54",  -- 84
        22588 => X"65",  -- 101
        22589 => X"75",  -- 117
        22590 => X"7E",  -- 126
        22591 => X"82",  -- 130
        22592 => X"87",  -- 135
        22593 => X"89",  -- 137
        22594 => X"8B",  -- 139
        22595 => X"8C",  -- 140
        22596 => X"8B",  -- 139
        22597 => X"91",  -- 145
        22598 => X"9E",  -- 158
        22599 => X"A8",  -- 168
        22600 => X"BA",  -- 186
        22601 => X"B2",  -- 178
        22602 => X"AC",  -- 172
        22603 => X"AC",  -- 172
        22604 => X"AF",  -- 175
        22605 => X"B2",  -- 178
        22606 => X"B4",  -- 180
        22607 => X"B7",  -- 183
        22608 => X"C1",  -- 193
        22609 => X"C4",  -- 196
        22610 => X"C9",  -- 201
        22611 => X"CC",  -- 204
        22612 => X"CD",  -- 205
        22613 => X"CD",  -- 205
        22614 => X"CD",  -- 205
        22615 => X"CE",  -- 206
        22616 => X"D0",  -- 208
        22617 => X"D2",  -- 210
        22618 => X"D0",  -- 208
        22619 => X"CA",  -- 202
        22620 => X"C3",  -- 195
        22621 => X"B8",  -- 184
        22622 => X"A5",  -- 165
        22623 => X"94",  -- 148
        22624 => X"86",  -- 134
        22625 => X"89",  -- 137
        22626 => X"8E",  -- 142
        22627 => X"97",  -- 151
        22628 => X"A4",  -- 164
        22629 => X"AE",  -- 174
        22630 => X"AE",  -- 174
        22631 => X"A7",  -- 167
        22632 => X"AA",  -- 170
        22633 => X"AA",  -- 170
        22634 => X"AA",  -- 170
        22635 => X"A7",  -- 167
        22636 => X"A4",  -- 164
        22637 => X"A1",  -- 161
        22638 => X"9F",  -- 159
        22639 => X"9E",  -- 158
        22640 => X"A2",  -- 162
        22641 => X"97",  -- 151
        22642 => X"90",  -- 144
        22643 => X"8B",  -- 139
        22644 => X"81",  -- 129
        22645 => X"75",  -- 117
        22646 => X"61",  -- 97
        22647 => X"46",  -- 70
        22648 => X"30",  -- 48
        22649 => X"39",  -- 57
        22650 => X"46",  -- 70
        22651 => X"56",  -- 86
        22652 => X"6A",  -- 106
        22653 => X"82",  -- 130
        22654 => X"93",  -- 147
        22655 => X"9B",  -- 155
        22656 => X"9B",  -- 155
        22657 => X"98",  -- 152
        22658 => X"95",  -- 149
        22659 => X"95",  -- 149
        22660 => X"98",  -- 152
        22661 => X"9D",  -- 157
        22662 => X"A4",  -- 164
        22663 => X"A8",  -- 168
        22664 => X"A9",  -- 169
        22665 => X"A9",  -- 169
        22666 => X"AA",  -- 170
        22667 => X"B0",  -- 176
        22668 => X"B9",  -- 185
        22669 => X"BD",  -- 189
        22670 => X"BB",  -- 187
        22671 => X"B9",  -- 185
        22672 => X"B8",  -- 184
        22673 => X"B7",  -- 183
        22674 => X"AB",  -- 171
        22675 => X"88",  -- 136
        22676 => X"52",  -- 82
        22677 => X"2C",  -- 44
        22678 => X"2E",  -- 46
        22679 => X"42",  -- 66
        22680 => X"6A",  -- 106
        22681 => X"7B",  -- 123
        22682 => X"88",  -- 136
        22683 => X"8B",  -- 139
        22684 => X"8B",  -- 139
        22685 => X"8C",  -- 140
        22686 => X"89",  -- 137
        22687 => X"84",  -- 132
        22688 => X"8E",  -- 142
        22689 => X"82",  -- 130
        22690 => X"7B",  -- 123
        22691 => X"80",  -- 128
        22692 => X"8A",  -- 138
        22693 => X"94",  -- 148
        22694 => X"9F",  -- 159
        22695 => X"AB",  -- 171
        22696 => X"AA",  -- 170
        22697 => X"A9",  -- 169
        22698 => X"AD",  -- 173
        22699 => X"B1",  -- 177
        22700 => X"B0",  -- 176
        22701 => X"A7",  -- 167
        22702 => X"9D",  -- 157
        22703 => X"96",  -- 150
        22704 => X"A3",  -- 163
        22705 => X"AD",  -- 173
        22706 => X"AF",  -- 175
        22707 => X"B0",  -- 176
        22708 => X"B7",  -- 183
        22709 => X"B4",  -- 180
        22710 => X"97",  -- 151
        22711 => X"71",  -- 113
        22712 => X"7A",  -- 122
        22713 => X"9E",  -- 158
        22714 => X"B1",  -- 177
        22715 => X"AA",  -- 170
        22716 => X"A0",  -- 160
        22717 => X"9F",  -- 159
        22718 => X"A7",  -- 167
        22719 => X"B3",  -- 179
        22720 => X"B0",  -- 176
        22721 => X"B2",  -- 178
        22722 => X"B2",  -- 178
        22723 => X"B2",  -- 178
        22724 => X"B0",  -- 176
        22725 => X"AC",  -- 172
        22726 => X"AA",  -- 170
        22727 => X"A7",  -- 167
        22728 => X"A7",  -- 167
        22729 => X"A3",  -- 163
        22730 => X"9D",  -- 157
        22731 => X"99",  -- 153
        22732 => X"99",  -- 153
        22733 => X"9A",  -- 154
        22734 => X"9B",  -- 155
        22735 => X"9A",  -- 154
        22736 => X"97",  -- 151
        22737 => X"89",  -- 137
        22738 => X"80",  -- 128
        22739 => X"82",  -- 130
        22740 => X"82",  -- 130
        22741 => X"7E",  -- 126
        22742 => X"7F",  -- 127
        22743 => X"86",  -- 134
        22744 => X"82",  -- 130
        22745 => X"87",  -- 135
        22746 => X"78",  -- 120
        22747 => X"6C",  -- 108
        22748 => X"67",  -- 103
        22749 => X"43",  -- 67
        22750 => X"22",  -- 34
        22751 => X"27",  -- 39
        22752 => X"45",  -- 69
        22753 => X"4E",  -- 78
        22754 => X"40",  -- 64
        22755 => X"2B",  -- 43
        22756 => X"23",  -- 35
        22757 => X"1D",  -- 29
        22758 => X"27",  -- 39
        22759 => X"42",  -- 66
        22760 => X"4A",  -- 74
        22761 => X"51",  -- 81
        22762 => X"52",  -- 82
        22763 => X"52",  -- 82
        22764 => X"4A",  -- 74
        22765 => X"3D",  -- 61
        22766 => X"42",  -- 66
        22767 => X"56",  -- 86
        22768 => X"61",  -- 97
        22769 => X"59",  -- 89
        22770 => X"4E",  -- 78
        22771 => X"5C",  -- 92
        22772 => X"84",  -- 132
        22773 => X"9E",  -- 158
        22774 => X"7F",  -- 127
        22775 => X"4B",  -- 75
        22776 => X"29",  -- 41
        22777 => X"1F",  -- 31
        22778 => X"18",  -- 24
        22779 => X"22",  -- 34
        22780 => X"5B",  -- 91
        22781 => X"65",  -- 101
        22782 => X"65",  -- 101
        22783 => X"67",  -- 103
        22784 => X"78",  -- 120
        22785 => X"78",  -- 120
        22786 => X"75",  -- 117
        22787 => X"69",  -- 105
        22788 => X"59",  -- 89
        22789 => X"4E",  -- 78
        22790 => X"51",  -- 81
        22791 => X"5B",  -- 91
        22792 => X"6F",  -- 111
        22793 => X"71",  -- 113
        22794 => X"95",  -- 149
        22795 => X"8B",  -- 139
        22796 => X"98",  -- 152
        22797 => X"96",  -- 150
        22798 => X"89",  -- 137
        22799 => X"86",  -- 134
        22800 => X"66",  -- 102
        22801 => X"5E",  -- 94
        22802 => X"59",  -- 89
        22803 => X"53",  -- 83
        22804 => X"44",  -- 68
        22805 => X"44",  -- 68
        22806 => X"66",  -- 102
        22807 => X"91",  -- 145
        22808 => X"92",  -- 146
        22809 => X"91",  -- 145
        22810 => X"79",  -- 121
        22811 => X"60",  -- 96
        22812 => X"38",  -- 56
        22813 => X"08",  -- 8
        22814 => X"23",  -- 35
        22815 => X"24",  -- 36
        22816 => X"28",  -- 40
        22817 => X"0F",  -- 15
        22818 => X"06",  -- 6
        22819 => X"11",  -- 17
        22820 => X"51",  -- 81
        22821 => X"78",  -- 120
        22822 => X"7F",  -- 127
        22823 => X"61",  -- 97
        22824 => X"38",  -- 56
        22825 => X"29",  -- 41
        22826 => X"0E",  -- 14
        22827 => X"12",  -- 18
        22828 => X"09",  -- 9
        22829 => X"11",  -- 17
        22830 => X"0B",  -- 11
        22831 => X"12",  -- 18
        22832 => X"27",  -- 39
        22833 => X"46",  -- 70
        22834 => X"62",  -- 98
        22835 => X"72",  -- 114
        22836 => X"84",  -- 132
        22837 => X"95",  -- 149
        22838 => X"8D",  -- 141
        22839 => X"79",  -- 121
        22840 => X"56",  -- 86
        22841 => X"3F",  -- 63
        22842 => X"45",  -- 69
        22843 => X"49",  -- 73
        22844 => X"2C",  -- 44
        22845 => X"28",  -- 40
        22846 => X"49",  -- 73
        22847 => X"60",  -- 96
        22848 => X"84",  -- 132
        22849 => X"7F",  -- 127
        22850 => X"89",  -- 137
        22851 => X"86",  -- 134
        22852 => X"56",  -- 86
        22853 => X"18",  -- 24
        22854 => X"09",  -- 9
        22855 => X"1E",  -- 30
        22856 => X"30",  -- 48
        22857 => X"3F",  -- 63
        22858 => X"50",  -- 80
        22859 => X"66",  -- 102
        22860 => X"83",  -- 131
        22861 => X"8E",  -- 142
        22862 => X"82",  -- 130
        22863 => X"79",  -- 121
        22864 => X"5D",  -- 93
        22865 => X"6B",  -- 107
        22866 => X"74",  -- 116
        22867 => X"7D",  -- 125
        22868 => X"63",  -- 99
        22869 => X"34",  -- 52
        22870 => X"1C",  -- 28
        22871 => X"0F",  -- 15
        22872 => X"13",  -- 19
        22873 => X"19",  -- 25
        22874 => X"35",  -- 53
        22875 => X"2B",  -- 43
        22876 => X"15",  -- 21
        22877 => X"1A",  -- 26
        22878 => X"24",  -- 36
        22879 => X"2A",  -- 42
        22880 => X"46",  -- 70
        22881 => X"5A",  -- 90
        22882 => X"7B",  -- 123
        22883 => X"82",  -- 130
        22884 => X"4E",  -- 78
        22885 => X"27",  -- 39
        22886 => X"5F",  -- 95
        22887 => X"A8",  -- 168
        22888 => X"9C",  -- 156
        22889 => X"A8",  -- 168
        22890 => X"97",  -- 151
        22891 => X"85",  -- 133
        22892 => X"84",  -- 132
        22893 => X"83",  -- 131
        22894 => X"8B",  -- 139
        22895 => X"A6",  -- 166
        22896 => X"92",  -- 146
        22897 => X"73",  -- 115
        22898 => X"59",  -- 89
        22899 => X"57",  -- 87
        22900 => X"5B",  -- 91
        22901 => X"52",  -- 82
        22902 => X"3F",  -- 63
        22903 => X"32",  -- 50
        22904 => X"22",  -- 34
        22905 => X"22",  -- 34
        22906 => X"24",  -- 36
        22907 => X"2E",  -- 46
        22908 => X"42",  -- 66
        22909 => X"5B",  -- 91
        22910 => X"75",  -- 117
        22911 => X"84",  -- 132
        22912 => X"86",  -- 134
        22913 => X"87",  -- 135
        22914 => X"86",  -- 134
        22915 => X"86",  -- 134
        22916 => X"89",  -- 137
        22917 => X"93",  -- 147
        22918 => X"9F",  -- 159
        22919 => X"A8",  -- 168
        22920 => X"B0",  -- 176
        22921 => X"AA",  -- 170
        22922 => X"A8",  -- 168
        22923 => X"AD",  -- 173
        22924 => X"B0",  -- 176
        22925 => X"B3",  -- 179
        22926 => X"B6",  -- 182
        22927 => X"B9",  -- 185
        22928 => X"BC",  -- 188
        22929 => X"BF",  -- 191
        22930 => X"C4",  -- 196
        22931 => X"C6",  -- 198
        22932 => X"C7",  -- 199
        22933 => X"C8",  -- 200
        22934 => X"C8",  -- 200
        22935 => X"CA",  -- 202
        22936 => X"CB",  -- 203
        22937 => X"CA",  -- 202
        22938 => X"C6",  -- 198
        22939 => X"C1",  -- 193
        22940 => X"BB",  -- 187
        22941 => X"B2",  -- 178
        22942 => X"A0",  -- 160
        22943 => X"8E",  -- 142
        22944 => X"83",  -- 131
        22945 => X"8A",  -- 138
        22946 => X"93",  -- 147
        22947 => X"9D",  -- 157
        22948 => X"AA",  -- 170
        22949 => X"B2",  -- 178
        22950 => X"AE",  -- 174
        22951 => X"A7",  -- 167
        22952 => X"A6",  -- 166
        22953 => X"A7",  -- 167
        22954 => X"A7",  -- 167
        22955 => X"A7",  -- 167
        22956 => X"A6",  -- 166
        22957 => X"A7",  -- 167
        22958 => X"A8",  -- 168
        22959 => X"AA",  -- 170
        22960 => X"99",  -- 153
        22961 => X"8D",  -- 141
        22962 => X"8A",  -- 138
        22963 => X"8B",  -- 139
        22964 => X"87",  -- 135
        22965 => X"7D",  -- 125
        22966 => X"63",  -- 99
        22967 => X"41",  -- 65
        22968 => X"34",  -- 52
        22969 => X"2F",  -- 47
        22970 => X"31",  -- 49
        22971 => X"42",  -- 66
        22972 => X"66",  -- 102
        22973 => X"87",  -- 135
        22974 => X"93",  -- 147
        22975 => X"91",  -- 145
        22976 => X"9B",  -- 155
        22977 => X"98",  -- 152
        22978 => X"97",  -- 151
        22979 => X"9D",  -- 157
        22980 => X"A5",  -- 165
        22981 => X"AA",  -- 170
        22982 => X"A6",  -- 166
        22983 => X"A2",  -- 162
        22984 => X"AF",  -- 175
        22985 => X"AD",  -- 173
        22986 => X"B0",  -- 176
        22987 => X"B7",  -- 183
        22988 => X"C0",  -- 192
        22989 => X"C4",  -- 196
        22990 => X"BF",  -- 191
        22991 => X"BB",  -- 187
        22992 => X"B7",  -- 183
        22993 => X"B5",  -- 181
        22994 => X"B1",  -- 177
        22995 => X"95",  -- 149
        22996 => X"51",  -- 81
        22997 => X"1D",  -- 29
        22998 => X"2F",  -- 47
        22999 => X"65",  -- 101
        23000 => X"7E",  -- 126
        23001 => X"85",  -- 133
        23002 => X"89",  -- 137
        23003 => X"85",  -- 133
        23004 => X"85",  -- 133
        23005 => X"8C",  -- 140
        23006 => X"90",  -- 144
        23007 => X"8F",  -- 143
        23008 => X"7C",  -- 124
        23009 => X"7C",  -- 124
        23010 => X"86",  -- 134
        23011 => X"94",  -- 148
        23012 => X"99",  -- 153
        23013 => X"97",  -- 151
        23014 => X"9E",  -- 158
        23015 => X"A9",  -- 169
        23016 => X"AB",  -- 171
        23017 => X"AB",  -- 171
        23018 => X"AE",  -- 174
        23019 => X"B1",  -- 177
        23020 => X"AF",  -- 175
        23021 => X"A8",  -- 168
        23022 => X"A5",  -- 165
        23023 => X"A3",  -- 163
        23024 => X"A5",  -- 165
        23025 => X"AE",  -- 174
        23026 => X"B0",  -- 176
        23027 => X"B1",  -- 177
        23028 => X"BB",  -- 187
        23029 => X"BB",  -- 187
        23030 => X"9C",  -- 156
        23031 => X"74",  -- 116
        23032 => X"7E",  -- 126
        23033 => X"A2",  -- 162
        23034 => X"B8",  -- 184
        23035 => X"B4",  -- 180
        23036 => X"A8",  -- 168
        23037 => X"9D",  -- 157
        23038 => X"9B",  -- 155
        23039 => X"A2",  -- 162
        23040 => X"AE",  -- 174
        23041 => X"B0",  -- 176
        23042 => X"B2",  -- 178
        23043 => X"B1",  -- 177
        23044 => X"AF",  -- 175
        23045 => X"AC",  -- 172
        23046 => X"A9",  -- 169
        23047 => X"A9",  -- 169
        23048 => X"A5",  -- 165
        23049 => X"9D",  -- 157
        23050 => X"97",  -- 151
        23051 => X"95",  -- 149
        23052 => X"91",  -- 145
        23053 => X"8B",  -- 139
        23054 => X"88",  -- 136
        23055 => X"87",  -- 135
        23056 => X"79",  -- 121
        23057 => X"73",  -- 115
        23058 => X"6B",  -- 107
        23059 => X"68",  -- 104
        23060 => X"69",  -- 105
        23061 => X"69",  -- 105
        23062 => X"65",  -- 101
        23063 => X"60",  -- 96
        23064 => X"67",  -- 103
        23065 => X"62",  -- 98
        23066 => X"5F",  -- 95
        23067 => X"5F",  -- 95
        23068 => X"5C",  -- 92
        23069 => X"4E",  -- 78
        23070 => X"3A",  -- 58
        23071 => X"2B",  -- 43
        23072 => X"4A",  -- 74
        23073 => X"48",  -- 72
        23074 => X"40",  -- 64
        23075 => X"33",  -- 51
        23076 => X"28",  -- 40
        23077 => X"2A",  -- 42
        23078 => X"34",  -- 52
        23079 => X"3E",  -- 62
        23080 => X"3A",  -- 58
        23081 => X"4A",  -- 74
        23082 => X"41",  -- 65
        23083 => X"2D",  -- 45
        23084 => X"39",  -- 57
        23085 => X"57",  -- 87
        23086 => X"65",  -- 101
        23087 => X"63",  -- 99
        23088 => X"51",  -- 81
        23089 => X"68",  -- 104
        23090 => X"84",  -- 132
        23091 => X"A2",  -- 162
        23092 => X"AB",  -- 171
        23093 => X"7D",  -- 125
        23094 => X"40",  -- 64
        23095 => X"2A",  -- 42
        23096 => X"1D",  -- 29
        23097 => X"18",  -- 24
        23098 => X"2A",  -- 42
        23099 => X"53",  -- 83
        23100 => X"66",  -- 102
        23101 => X"5E",  -- 94
        23102 => X"5B",  -- 91
        23103 => X"65",  -- 101
        23104 => X"70",  -- 112
        23105 => X"5E",  -- 94
        23106 => X"71",  -- 113
        23107 => X"81",  -- 129
        23108 => X"73",  -- 115
        23109 => X"8A",  -- 138
        23110 => X"82",  -- 130
        23111 => X"88",  -- 136
        23112 => X"98",  -- 152
        23113 => X"A5",  -- 165
        23114 => X"9B",  -- 155
        23115 => X"8C",  -- 140
        23116 => X"62",  -- 98
        23117 => X"55",  -- 85
        23118 => X"3B",  -- 59
        23119 => X"30",  -- 48
        23120 => X"1E",  -- 30
        23121 => X"19",  -- 25
        23122 => X"1B",  -- 27
        23123 => X"1C",  -- 28
        23124 => X"18",  -- 24
        23125 => X"1C",  -- 28
        23126 => X"41",  -- 65
        23127 => X"6B",  -- 107
        23128 => X"79",  -- 121
        23129 => X"8C",  -- 140
        23130 => X"7E",  -- 126
        23131 => X"55",  -- 85
        23132 => X"0E",  -- 14
        23133 => X"19",  -- 25
        23134 => X"39",  -- 57
        23135 => X"1E",  -- 30
        23136 => X"30",  -- 48
        23137 => X"0D",  -- 13
        23138 => X"0F",  -- 15
        23139 => X"07",  -- 7
        23140 => X"21",  -- 33
        23141 => X"6B",  -- 107
        23142 => X"7E",  -- 126
        23143 => X"86",  -- 134
        23144 => X"6F",  -- 111
        23145 => X"3B",  -- 59
        23146 => X"14",  -- 20
        23147 => X"0C",  -- 12
        23148 => X"08",  -- 8
        23149 => X"04",  -- 4
        23150 => X"06",  -- 6
        23151 => X"09",  -- 9
        23152 => X"08",  -- 8
        23153 => X"12",  -- 18
        23154 => X"14",  -- 20
        23155 => X"3A",  -- 58
        23156 => X"5A",  -- 90
        23157 => X"6D",  -- 109
        23158 => X"8F",  -- 143
        23159 => X"97",  -- 151
        23160 => X"9D",  -- 157
        23161 => X"86",  -- 134
        23162 => X"87",  -- 135
        23163 => X"7D",  -- 125
        23164 => X"5A",  -- 90
        23165 => X"6E",  -- 110
        23166 => X"69",  -- 105
        23167 => X"6F",  -- 111
        23168 => X"7E",  -- 126
        23169 => X"87",  -- 135
        23170 => X"83",  -- 131
        23171 => X"6E",  -- 110
        23172 => X"5D",  -- 93
        23173 => X"35",  -- 53
        23174 => X"0B",  -- 11
        23175 => X"10",  -- 16
        23176 => X"1F",  -- 31
        23177 => X"24",  -- 36
        23178 => X"29",  -- 41
        23179 => X"38",  -- 56
        23180 => X"50",  -- 80
        23181 => X"61",  -- 97
        23182 => X"78",  -- 120
        23183 => X"92",  -- 146
        23184 => X"A0",  -- 160
        23185 => X"8C",  -- 140
        23186 => X"86",  -- 134
        23187 => X"93",  -- 147
        23188 => X"93",  -- 147
        23189 => X"79",  -- 121
        23190 => X"5A",  -- 90
        23191 => X"4C",  -- 76
        23192 => X"47",  -- 71
        23193 => X"34",  -- 52
        23194 => X"20",  -- 32
        23195 => X"1B",  -- 27
        23196 => X"1D",  -- 29
        23197 => X"25",  -- 37
        23198 => X"37",  -- 55
        23199 => X"49",  -- 73
        23200 => X"4B",  -- 75
        23201 => X"6E",  -- 110
        23202 => X"7C",  -- 124
        23203 => X"8E",  -- 142
        23204 => X"65",  -- 101
        23205 => X"38",  -- 56
        23206 => X"62",  -- 98
        23207 => X"8B",  -- 139
        23208 => X"98",  -- 152
        23209 => X"98",  -- 152
        23210 => X"8E",  -- 142
        23211 => X"7F",  -- 127
        23212 => X"7F",  -- 127
        23213 => X"89",  -- 137
        23214 => X"86",  -- 134
        23215 => X"79",  -- 121
        23216 => X"91",  -- 145
        23217 => X"7E",  -- 126
        23218 => X"63",  -- 99
        23219 => X"4E",  -- 78
        23220 => X"46",  -- 70
        23221 => X"42",  -- 66
        23222 => X"39",  -- 57
        23223 => X"30",  -- 48
        23224 => X"2E",  -- 46
        23225 => X"30",  -- 48
        23226 => X"27",  -- 39
        23227 => X"1D",  -- 29
        23228 => X"2A",  -- 42
        23229 => X"50",  -- 80
        23230 => X"73",  -- 115
        23231 => X"80",  -- 128
        23232 => X"82",  -- 130
        23233 => X"94",  -- 148
        23234 => X"9A",  -- 154
        23235 => X"91",  -- 145
        23236 => X"93",  -- 147
        23237 => X"A3",  -- 163
        23238 => X"AC",  -- 172
        23239 => X"AA",  -- 170
        23240 => X"B4",  -- 180
        23241 => X"B8",  -- 184
        23242 => X"BB",  -- 187
        23243 => X"B9",  -- 185
        23244 => X"B7",  -- 183
        23245 => X"B6",  -- 182
        23246 => X"BB",  -- 187
        23247 => X"BF",  -- 191
        23248 => X"C2",  -- 194
        23249 => X"C9",  -- 201
        23250 => X"D0",  -- 208
        23251 => X"D3",  -- 211
        23252 => X"D2",  -- 210
        23253 => X"D0",  -- 208
        23254 => X"CF",  -- 207
        23255 => X"D1",  -- 209
        23256 => X"CE",  -- 206
        23257 => X"D1",  -- 209
        23258 => X"D3",  -- 211
        23259 => X"CE",  -- 206
        23260 => X"C7",  -- 199
        23261 => X"BF",  -- 191
        23262 => X"B3",  -- 179
        23263 => X"AC",  -- 172
        23264 => X"9D",  -- 157
        23265 => X"90",  -- 144
        23266 => X"94",  -- 148
        23267 => X"A9",  -- 169
        23268 => X"BB",  -- 187
        23269 => X"B8",  -- 184
        23270 => X"AF",  -- 175
        23271 => X"AE",  -- 174
        23272 => X"A8",  -- 168
        23273 => X"A6",  -- 166
        23274 => X"A7",  -- 167
        23275 => X"AF",  -- 175
        23276 => X"B3",  -- 179
        23277 => X"AD",  -- 173
        23278 => X"A2",  -- 162
        23279 => X"9B",  -- 155
        23280 => X"8E",  -- 142
        23281 => X"8F",  -- 143
        23282 => X"8F",  -- 143
        23283 => X"8E",  -- 142
        23284 => X"8E",  -- 142
        23285 => X"82",  -- 130
        23286 => X"6C",  -- 108
        23287 => X"57",  -- 87
        23288 => X"3F",  -- 63
        23289 => X"33",  -- 51
        23290 => X"35",  -- 53
        23291 => X"50",  -- 80
        23292 => X"73",  -- 115
        23293 => X"89",  -- 137
        23294 => X"96",  -- 150
        23295 => X"9F",  -- 159
        23296 => X"9E",  -- 158
        23297 => X"A2",  -- 162
        23298 => X"A5",  -- 165
        23299 => X"A7",  -- 167
        23300 => X"A7",  -- 167
        23301 => X"A8",  -- 168
        23302 => X"AD",  -- 173
        23303 => X"AF",  -- 175
        23304 => X"B5",  -- 181
        23305 => X"B1",  -- 177
        23306 => X"B3",  -- 179
        23307 => X"BB",  -- 187
        23308 => X"C1",  -- 193
        23309 => X"C0",  -- 192
        23310 => X"BE",  -- 190
        23311 => X"BF",  -- 191
        23312 => X"C3",  -- 195
        23313 => X"B6",  -- 182
        23314 => X"A4",  -- 164
        23315 => X"72",  -- 114
        23316 => X"32",  -- 50
        23317 => X"31",  -- 49
        23318 => X"54",  -- 84
        23319 => X"65",  -- 101
        23320 => X"8A",  -- 138
        23321 => X"89",  -- 137
        23322 => X"8A",  -- 138
        23323 => X"8F",  -- 143
        23324 => X"96",  -- 150
        23325 => X"96",  -- 150
        23326 => X"8D",  -- 141
        23327 => X"83",  -- 131
        23328 => X"89",  -- 137
        23329 => X"89",  -- 137
        23330 => X"8B",  -- 139
        23331 => X"95",  -- 149
        23332 => X"9A",  -- 154
        23333 => X"97",  -- 151
        23334 => X"9E",  -- 158
        23335 => X"B2",  -- 178
        23336 => X"B4",  -- 180
        23337 => X"AB",  -- 171
        23338 => X"A7",  -- 167
        23339 => X"AD",  -- 173
        23340 => X"AF",  -- 175
        23341 => X"AA",  -- 170
        23342 => X"A1",  -- 161
        23343 => X"9D",  -- 157
        23344 => X"AF",  -- 175
        23345 => X"AF",  -- 175
        23346 => X"B2",  -- 178
        23347 => X"B9",  -- 185
        23348 => X"BF",  -- 191
        23349 => X"B1",  -- 177
        23350 => X"8E",  -- 142
        23351 => X"6F",  -- 111
        23352 => X"7C",  -- 124
        23353 => X"98",  -- 152
        23354 => X"B1",  -- 177
        23355 => X"B2",  -- 178
        23356 => X"AD",  -- 173
        23357 => X"AA",  -- 170
        23358 => X"A6",  -- 166
        23359 => X"A2",  -- 162
        23360 => X"AD",  -- 173
        23361 => X"AE",  -- 174
        23362 => X"AF",  -- 175
        23363 => X"AE",  -- 174
        23364 => X"AB",  -- 171
        23365 => X"A6",  -- 166
        23366 => X"A3",  -- 163
        23367 => X"A1",  -- 161
        23368 => X"A2",  -- 162
        23369 => X"9C",  -- 156
        23370 => X"97",  -- 151
        23371 => X"95",  -- 149
        23372 => X"8F",  -- 143
        23373 => X"85",  -- 133
        23374 => X"7E",  -- 126
        23375 => X"7C",  -- 124
        23376 => X"6D",  -- 109
        23377 => X"66",  -- 102
        23378 => X"60",  -- 96
        23379 => X"5E",  -- 94
        23380 => X"5F",  -- 95
        23381 => X"5E",  -- 94
        23382 => X"59",  -- 89
        23383 => X"55",  -- 85
        23384 => X"52",  -- 82
        23385 => X"52",  -- 82
        23386 => X"55",  -- 85
        23387 => X"5B",  -- 91
        23388 => X"5A",  -- 90
        23389 => X"53",  -- 83
        23390 => X"4B",  -- 75
        23391 => X"48",  -- 72
        23392 => X"59",  -- 89
        23393 => X"55",  -- 85
        23394 => X"4A",  -- 74
        23395 => X"3B",  -- 59
        23396 => X"32",  -- 50
        23397 => X"31",  -- 49
        23398 => X"32",  -- 50
        23399 => X"30",  -- 48
        23400 => X"45",  -- 69
        23401 => X"3C",  -- 60
        23402 => X"35",  -- 53
        23403 => X"46",  -- 70
        23404 => X"65",  -- 101
        23405 => X"6B",  -- 107
        23406 => X"53",  -- 83
        23407 => X"42",  -- 66
        23408 => X"4A",  -- 74
        23409 => X"7C",  -- 124
        23410 => X"A2",  -- 162
        23411 => X"A2",  -- 162
        23412 => X"89",  -- 137
        23413 => X"5B",  -- 91
        23414 => X"33",  -- 51
        23415 => X"2A",  -- 42
        23416 => X"27",  -- 39
        23417 => X"3E",  -- 62
        23418 => X"58",  -- 88
        23419 => X"5F",  -- 95
        23420 => X"53",  -- 83
        23421 => X"4E",  -- 78
        23422 => X"63",  -- 99
        23423 => X"7E",  -- 126
        23424 => X"73",  -- 115
        23425 => X"68",  -- 104
        23426 => X"6D",  -- 109
        23427 => X"80",  -- 128
        23428 => X"8F",  -- 143
        23429 => X"A0",  -- 160
        23430 => X"9B",  -- 155
        23431 => X"A1",  -- 161
        23432 => X"C3",  -- 195
        23433 => X"A7",  -- 167
        23434 => X"76",  -- 118
        23435 => X"49",  -- 73
        23436 => X"22",  -- 34
        23437 => X"16",  -- 22
        23438 => X"09",  -- 9
        23439 => X"04",  -- 4
        23440 => X"06",  -- 6
        23441 => X"03",  -- 3
        23442 => X"09",  -- 9
        23443 => X"15",  -- 21
        23444 => X"19",  -- 25
        23445 => X"19",  -- 25
        23446 => X"24",  -- 36
        23447 => X"35",  -- 53
        23448 => X"59",  -- 89
        23449 => X"82",  -- 130
        23450 => X"70",  -- 112
        23451 => X"43",  -- 67
        23452 => X"0D",  -- 13
        23453 => X"17",  -- 23
        23454 => X"2F",  -- 47
        23455 => X"25",  -- 37
        23456 => X"49",  -- 73
        23457 => X"04",  -- 4
        23458 => X"0C",  -- 12
        23459 => X"12",  -- 18
        23460 => X"0B",  -- 11
        23461 => X"3D",  -- 61
        23462 => X"7F",  -- 127
        23463 => X"99",  -- 153
        23464 => X"89",  -- 137
        23465 => X"54",  -- 84
        23466 => X"22",  -- 34
        23467 => X"0F",  -- 15
        23468 => X"0B",  -- 11
        23469 => X"0E",  -- 14
        23470 => X"0B",  -- 11
        23471 => X"00",  -- 0
        23472 => X"04",  -- 4
        23473 => X"0D",  -- 13
        23474 => X"03",  -- 3
        23475 => X"03",  -- 3
        23476 => X"0D",  -- 13
        23477 => X"46",  -- 70
        23478 => X"8C",  -- 140
        23479 => X"AB",  -- 171
        23480 => X"B0",  -- 176
        23481 => X"A2",  -- 162
        23482 => X"96",  -- 150
        23483 => X"96",  -- 150
        23484 => X"89",  -- 137
        23485 => X"92",  -- 146
        23486 => X"80",  -- 128
        23487 => X"7B",  -- 123
        23488 => X"81",  -- 129
        23489 => X"66",  -- 102
        23490 => X"71",  -- 113
        23491 => X"78",  -- 120
        23492 => X"6A",  -- 106
        23493 => X"58",  -- 88
        23494 => X"2C",  -- 44
        23495 => X"07",  -- 7
        23496 => X"06",  -- 6
        23497 => X"13",  -- 19
        23498 => X"23",  -- 35
        23499 => X"33",  -- 51
        23500 => X"3E",  -- 62
        23501 => X"45",  -- 69
        23502 => X"5E",  -- 94
        23503 => X"80",  -- 128
        23504 => X"97",  -- 151
        23505 => X"8D",  -- 141
        23506 => X"85",  -- 133
        23507 => X"84",  -- 132
        23508 => X"89",  -- 137
        23509 => X"8E",  -- 142
        23510 => X"90",  -- 144
        23511 => X"8E",  -- 142
        23512 => X"5C",  -- 92
        23513 => X"4C",  -- 76
        23514 => X"33",  -- 51
        23515 => X"1E",  -- 30
        23516 => X"1D",  -- 29
        23517 => X"36",  -- 54
        23518 => X"57",  -- 87
        23519 => X"6F",  -- 111
        23520 => X"68",  -- 104
        23521 => X"79",  -- 121
        23522 => X"88",  -- 136
        23523 => X"A8",  -- 168
        23524 => X"8A",  -- 138
        23525 => X"57",  -- 87
        23526 => X"65",  -- 101
        23527 => X"70",  -- 112
        23528 => X"88",  -- 136
        23529 => X"97",  -- 151
        23530 => X"9D",  -- 157
        23531 => X"8E",  -- 142
        23532 => X"81",  -- 129
        23533 => X"83",  -- 131
        23534 => X"86",  -- 134
        23535 => X"85",  -- 133
        23536 => X"76",  -- 118
        23537 => X"70",  -- 112
        23538 => X"66",  -- 102
        23539 => X"5C",  -- 92
        23540 => X"54",  -- 84
        23541 => X"47",  -- 71
        23542 => X"34",  -- 52
        23543 => X"23",  -- 35
        23544 => X"26",  -- 38
        23545 => X"2A",  -- 42
        23546 => X"22",  -- 34
        23547 => X"19",  -- 25
        23548 => X"1F",  -- 31
        23549 => X"39",  -- 57
        23550 => X"59",  -- 89
        23551 => X"6A",  -- 106
        23552 => X"6D",  -- 109
        23553 => X"83",  -- 131
        23554 => X"94",  -- 148
        23555 => X"98",  -- 152
        23556 => X"9B",  -- 155
        23557 => X"A6",  -- 166
        23558 => X"AE",  -- 174
        23559 => X"AD",  -- 173
        23560 => X"B7",  -- 183
        23561 => X"B8",  -- 184
        23562 => X"BA",  -- 186
        23563 => X"BB",  -- 187
        23564 => X"BB",  -- 187
        23565 => X"BD",  -- 189
        23566 => X"C1",  -- 193
        23567 => X"C5",  -- 197
        23568 => X"C5",  -- 197
        23569 => X"C9",  -- 201
        23570 => X"CE",  -- 206
        23571 => X"CE",  -- 206
        23572 => X"CC",  -- 204
        23573 => X"C9",  -- 201
        23574 => X"CA",  -- 202
        23575 => X"CD",  -- 205
        23576 => X"CB",  -- 203
        23577 => X"CC",  -- 204
        23578 => X"CE",  -- 206
        23579 => X"CD",  -- 205
        23580 => X"CD",  -- 205
        23581 => X"C9",  -- 201
        23582 => X"BE",  -- 190
        23583 => X"B2",  -- 178
        23584 => X"95",  -- 149
        23585 => X"8A",  -- 138
        23586 => X"8A",  -- 138
        23587 => X"A0",  -- 160
        23588 => X"AF",  -- 175
        23589 => X"AE",  -- 174
        23590 => X"A8",  -- 168
        23591 => X"A5",  -- 165
        23592 => X"A7",  -- 167
        23593 => X"A6",  -- 166
        23594 => X"A5",  -- 165
        23595 => X"A5",  -- 165
        23596 => X"A8",  -- 168
        23597 => X"AA",  -- 170
        23598 => X"AA",  -- 170
        23599 => X"AA",  -- 170
        23600 => X"AD",  -- 173
        23601 => X"9F",  -- 159
        23602 => X"93",  -- 147
        23603 => X"91",  -- 145
        23604 => X"97",  -- 151
        23605 => X"90",  -- 144
        23606 => X"71",  -- 113
        23607 => X"52",  -- 82
        23608 => X"41",  -- 65
        23609 => X"34",  -- 52
        23610 => X"36",  -- 54
        23611 => X"50",  -- 80
        23612 => X"6F",  -- 111
        23613 => X"84",  -- 132
        23614 => X"8B",  -- 139
        23615 => X"8E",  -- 142
        23616 => X"9A",  -- 154
        23617 => X"9F",  -- 159
        23618 => X"A5",  -- 165
        23619 => X"A7",  -- 167
        23620 => X"AA",  -- 170
        23621 => X"AB",  -- 171
        23622 => X"AE",  -- 174
        23623 => X"B1",  -- 177
        23624 => X"B2",  -- 178
        23625 => X"B1",  -- 177
        23626 => X"B6",  -- 182
        23627 => X"C0",  -- 192
        23628 => X"C5",  -- 197
        23629 => X"C4",  -- 196
        23630 => X"C2",  -- 194
        23631 => X"C3",  -- 195
        23632 => X"B9",  -- 185
        23633 => X"B0",  -- 176
        23634 => X"9E",  -- 158
        23635 => X"73",  -- 115
        23636 => X"3E",  -- 62
        23637 => X"3C",  -- 60
        23638 => X"60",  -- 96
        23639 => X"78",  -- 120
        23640 => X"86",  -- 134
        23641 => X"88",  -- 136
        23642 => X"8F",  -- 143
        23643 => X"94",  -- 148
        23644 => X"98",  -- 152
        23645 => X"95",  -- 149
        23646 => X"8E",  -- 142
        23647 => X"87",  -- 135
        23648 => X"8E",  -- 142
        23649 => X"96",  -- 150
        23650 => X"96",  -- 150
        23651 => X"94",  -- 148
        23652 => X"98",  -- 152
        23653 => X"97",  -- 151
        23654 => X"99",  -- 153
        23655 => X"A5",  -- 165
        23656 => X"B2",  -- 178
        23657 => X"AC",  -- 172
        23658 => X"A9",  -- 169
        23659 => X"A9",  -- 169
        23660 => X"A6",  -- 166
        23661 => X"A3",  -- 163
        23662 => X"A3",  -- 163
        23663 => X"A8",  -- 168
        23664 => X"AF",  -- 175
        23665 => X"AE",  -- 174
        23666 => X"B1",  -- 177
        23667 => X"B9",  -- 185
        23668 => X"BF",  -- 191
        23669 => X"B6",  -- 182
        23670 => X"99",  -- 153
        23671 => X"7D",  -- 125
        23672 => X"8C",  -- 140
        23673 => X"9E",  -- 158
        23674 => X"AA",  -- 170
        23675 => X"AB",  -- 171
        23676 => X"AA",  -- 170
        23677 => X"AC",  -- 172
        23678 => X"AC",  -- 172
        23679 => X"A8",  -- 168
        23680 => X"AB",  -- 171
        23681 => X"AB",  -- 171
        23682 => X"AB",  -- 171
        23683 => X"A8",  -- 168
        23684 => X"A2",  -- 162
        23685 => X"9B",  -- 155
        23686 => X"96",  -- 150
        23687 => X"92",  -- 146
        23688 => X"94",  -- 148
        23689 => X"90",  -- 144
        23690 => X"8C",  -- 140
        23691 => X"8C",  -- 140
        23692 => X"88",  -- 136
        23693 => X"7E",  -- 126
        23694 => X"75",  -- 117
        23695 => X"70",  -- 112
        23696 => X"68",  -- 104
        23697 => X"63",  -- 99
        23698 => X"5D",  -- 93
        23699 => X"5B",  -- 91
        23700 => X"5D",  -- 93
        23701 => X"5D",  -- 93
        23702 => X"58",  -- 88
        23703 => X"55",  -- 85
        23704 => X"50",  -- 80
        23705 => X"52",  -- 82
        23706 => X"58",  -- 88
        23707 => X"5A",  -- 90
        23708 => X"57",  -- 87
        23709 => X"53",  -- 83
        23710 => X"52",  -- 82
        23711 => X"56",  -- 86
        23712 => X"67",  -- 103
        23713 => X"64",  -- 100
        23714 => X"56",  -- 86
        23715 => X"44",  -- 68
        23716 => X"3B",  -- 59
        23717 => X"3A",  -- 58
        23718 => X"33",  -- 51
        23719 => X"27",  -- 39
        23720 => X"16",  -- 22
        23721 => X"1A",  -- 26
        23722 => X"2D",  -- 45
        23723 => X"4B",  -- 75
        23724 => X"57",  -- 87
        23725 => X"47",  -- 71
        23726 => X"44",  -- 68
        23727 => X"5A",  -- 90
        23728 => X"70",  -- 112
        23729 => X"80",  -- 128
        23730 => X"84",  -- 132
        23731 => X"73",  -- 115
        23732 => X"5A",  -- 90
        23733 => X"3D",  -- 61
        23734 => X"2F",  -- 47
        23735 => X"33",  -- 51
        23736 => X"46",  -- 70
        23737 => X"58",  -- 88
        23738 => X"5B",  -- 91
        23739 => X"43",  -- 67
        23740 => X"3A",  -- 58
        23741 => X"4F",  -- 79
        23742 => X"6F",  -- 111
        23743 => X"82",  -- 130
        23744 => X"77",  -- 119
        23745 => X"7D",  -- 125
        23746 => X"7C",  -- 124
        23747 => X"8B",  -- 139
        23748 => X"AC",  -- 172
        23749 => X"B2",  -- 178
        23750 => X"B6",  -- 182
        23751 => X"AF",  -- 175
        23752 => X"B4",  -- 180
        23753 => X"7F",  -- 127
        23754 => X"42",  -- 66
        23755 => X"12",  -- 18
        23756 => X"06",  -- 6
        23757 => X"05",  -- 5
        23758 => X"07",  -- 7
        23759 => X"05",  -- 5
        23760 => X"06",  -- 6
        23761 => X"02",  -- 2
        23762 => X"01",  -- 1
        23763 => X"03",  -- 3
        23764 => X"09",  -- 9
        23765 => X"0E",  -- 14
        23766 => X"15",  -- 21
        23767 => X"19",  -- 25
        23768 => X"37",  -- 55
        23769 => X"69",  -- 105
        23770 => X"51",  -- 81
        23771 => X"23",  -- 35
        23772 => X"09",  -- 9
        23773 => X"1D",  -- 29
        23774 => X"2F",  -- 47
        23775 => X"35",  -- 53
        23776 => X"45",  -- 69
        23777 => X"0D",  -- 13
        23778 => X"12",  -- 18
        23779 => X"06",  -- 6
        23780 => X"09",  -- 9
        23781 => X"17",  -- 23
        23782 => X"4A",  -- 74
        23783 => X"78",  -- 120
        23784 => X"82",  -- 130
        23785 => X"77",  -- 119
        23786 => X"61",  -- 97
        23787 => X"3B",  -- 59
        23788 => X"14",  -- 20
        23789 => X"06",  -- 6
        23790 => X"0A",  -- 10
        23791 => X"0A",  -- 10
        23792 => X"08",  -- 8
        23793 => X"07",  -- 7
        23794 => X"0D",  -- 13
        23795 => X"07",  -- 7
        23796 => X"03",  -- 3
        23797 => X"14",  -- 20
        23798 => X"3D",  -- 61
        23799 => X"6D",  -- 109
        23800 => X"A7",  -- 167
        23801 => X"C0",  -- 192
        23802 => X"B1",  -- 177
        23803 => X"AE",  -- 174
        23804 => X"AD",  -- 173
        23805 => X"A3",  -- 163
        23806 => X"89",  -- 137
        23807 => X"7F",  -- 127
        23808 => X"7F",  -- 127
        23809 => X"83",  -- 131
        23810 => X"92",  -- 146
        23811 => X"75",  -- 117
        23812 => X"51",  -- 81
        23813 => X"53",  -- 83
        23814 => X"41",  -- 65
        23815 => X"1E",  -- 30
        23816 => X"0D",  -- 13
        23817 => X"18",  -- 24
        23818 => X"22",  -- 34
        23819 => X"29",  -- 41
        23820 => X"29",  -- 41
        23821 => X"22",  -- 34
        23822 => X"30",  -- 48
        23823 => X"4D",  -- 77
        23824 => X"5E",  -- 94
        23825 => X"77",  -- 119
        23826 => X"8E",  -- 142
        23827 => X"90",  -- 144
        23828 => X"8C",  -- 140
        23829 => X"84",  -- 132
        23830 => X"71",  -- 113
        23831 => X"5B",  -- 91
        23832 => X"6F",  -- 111
        23833 => X"6C",  -- 108
        23834 => X"55",  -- 85
        23835 => X"36",  -- 54
        23836 => X"26",  -- 38
        23837 => X"31",  -- 49
        23838 => X"47",  -- 71
        23839 => X"54",  -- 84
        23840 => X"6F",  -- 111
        23841 => X"81",  -- 129
        23842 => X"98",  -- 152
        23843 => X"B2",  -- 178
        23844 => X"8E",  -- 142
        23845 => X"60",  -- 96
        23846 => X"6F",  -- 111
        23847 => X"72",  -- 114
        23848 => X"7C",  -- 124
        23849 => X"95",  -- 149
        23850 => X"A5",  -- 165
        23851 => X"9D",  -- 157
        23852 => X"8C",  -- 140
        23853 => X"88",  -- 136
        23854 => X"8D",  -- 141
        23855 => X"90",  -- 144
        23856 => X"7E",  -- 126
        23857 => X"7C",  -- 124
        23858 => X"74",  -- 116
        23859 => X"69",  -- 105
        23860 => X"5C",  -- 92
        23861 => X"50",  -- 80
        23862 => X"3E",  -- 62
        23863 => X"2F",  -- 47
        23864 => X"2D",  -- 45
        23865 => X"2D",  -- 45
        23866 => X"27",  -- 39
        23867 => X"22",  -- 34
        23868 => X"23",  -- 35
        23869 => X"30",  -- 48
        23870 => X"4E",  -- 78
        23871 => X"68",  -- 104
        23872 => X"72",  -- 114
        23873 => X"7F",  -- 127
        23874 => X"8B",  -- 139
        23875 => X"91",  -- 145
        23876 => X"95",  -- 149
        23877 => X"9F",  -- 159
        23878 => X"AB",  -- 171
        23879 => X"B4",  -- 180
        23880 => X"B2",  -- 178
        23881 => X"B3",  -- 179
        23882 => X"B5",  -- 181
        23883 => X"B7",  -- 183
        23884 => X"BA",  -- 186
        23885 => X"BE",  -- 190
        23886 => X"C1",  -- 193
        23887 => X"C3",  -- 195
        23888 => X"BE",  -- 190
        23889 => X"C1",  -- 193
        23890 => X"C5",  -- 197
        23891 => X"C7",  -- 199
        23892 => X"C8",  -- 200
        23893 => X"CA",  -- 202
        23894 => X"CC",  -- 204
        23895 => X"D0",  -- 208
        23896 => X"D1",  -- 209
        23897 => X"D1",  -- 209
        23898 => X"CF",  -- 207
        23899 => X"CF",  -- 207
        23900 => X"CF",  -- 207
        23901 => X"CB",  -- 203
        23902 => X"BC",  -- 188
        23903 => X"AF",  -- 175
        23904 => X"93",  -- 147
        23905 => X"89",  -- 137
        23906 => X"89",  -- 137
        23907 => X"9D",  -- 157
        23908 => X"AC",  -- 172
        23909 => X"AE",  -- 174
        23910 => X"A9",  -- 169
        23911 => X"A7",  -- 167
        23912 => X"A1",  -- 161
        23913 => X"A8",  -- 168
        23914 => X"AC",  -- 172
        23915 => X"A9",  -- 169
        23916 => X"A7",  -- 167
        23917 => X"A9",  -- 169
        23918 => X"A6",  -- 166
        23919 => X"A0",  -- 160
        23920 => X"96",  -- 150
        23921 => X"95",  -- 149
        23922 => X"95",  -- 149
        23923 => X"98",  -- 152
        23924 => X"9A",  -- 154
        23925 => X"90",  -- 144
        23926 => X"7A",  -- 122
        23927 => X"64",  -- 100
        23928 => X"4C",  -- 76
        23929 => X"42",  -- 66
        23930 => X"42",  -- 66
        23931 => X"59",  -- 89
        23932 => X"79",  -- 121
        23933 => X"8C",  -- 140
        23934 => X"92",  -- 146
        23935 => X"93",  -- 147
        23936 => X"98",  -- 152
        23937 => X"9E",  -- 158
        23938 => X"A5",  -- 165
        23939 => X"AA",  -- 170
        23940 => X"AC",  -- 172
        23941 => X"AF",  -- 175
        23942 => X"B1",  -- 177
        23943 => X"B4",  -- 180
        23944 => X"B4",  -- 180
        23945 => X"B7",  -- 183
        23946 => X"BF",  -- 191
        23947 => X"C6",  -- 198
        23948 => X"C7",  -- 199
        23949 => X"C4",  -- 196
        23950 => X"C3",  -- 195
        23951 => X"C4",  -- 196
        23952 => X"BF",  -- 191
        23953 => X"B7",  -- 183
        23954 => X"8E",  -- 142
        23955 => X"52",  -- 82
        23956 => X"30",  -- 48
        23957 => X"43",  -- 67
        23958 => X"6D",  -- 109
        23959 => X"84",  -- 132
        23960 => X"92",  -- 146
        23961 => X"94",  -- 148
        23962 => X"97",  -- 151
        23963 => X"98",  -- 152
        23964 => X"97",  -- 151
        23965 => X"97",  -- 151
        23966 => X"99",  -- 153
        23967 => X"9B",  -- 155
        23968 => X"9C",  -- 156
        23969 => X"AB",  -- 171
        23970 => X"AF",  -- 175
        23971 => X"AB",  -- 171
        23972 => X"AE",  -- 174
        23973 => X"AD",  -- 173
        23974 => X"AA",  -- 170
        23975 => X"AC",  -- 172
        23976 => X"B8",  -- 184
        23977 => X"B7",  -- 183
        23978 => X"B4",  -- 180
        23979 => X"AD",  -- 173
        23980 => X"A2",  -- 162
        23981 => X"9C",  -- 156
        23982 => X"A1",  -- 161
        23983 => X"A7",  -- 167
        23984 => X"AE",  -- 174
        23985 => X"AE",  -- 174
        23986 => X"B2",  -- 178
        23987 => X"B9",  -- 185
        23988 => X"C1",  -- 193
        23989 => X"BE",  -- 190
        23990 => X"A8",  -- 168
        23991 => X"93",  -- 147
        23992 => X"9D",  -- 157
        23993 => X"A1",  -- 161
        23994 => X"A1",  -- 161
        23995 => X"A0",  -- 160
        23996 => X"A3",  -- 163
        23997 => X"AC",  -- 172
        23998 => X"AF",  -- 175
        23999 => X"AC",  -- 172
        24000 => X"A3",  -- 163
        24001 => X"A5",  -- 165
        24002 => X"A5",  -- 165
        24003 => X"A2",  -- 162
        24004 => X"99",  -- 153
        24005 => X"8D",  -- 141
        24006 => X"84",  -- 132
        24007 => X"7D",  -- 125
        24008 => X"7B",  -- 123
        24009 => X"76",  -- 118
        24010 => X"75",  -- 117
        24011 => X"79",  -- 121
        24012 => X"79",  -- 121
        24013 => X"73",  -- 115
        24014 => X"6C",  -- 108
        24015 => X"69",  -- 105
        24016 => X"69",  -- 105
        24017 => X"65",  -- 101
        24018 => X"60",  -- 96
        24019 => X"5E",  -- 94
        24020 => X"60",  -- 96
        24021 => X"5F",  -- 95
        24022 => X"5C",  -- 92
        24023 => X"5A",  -- 90
        24024 => X"59",  -- 89
        24025 => X"59",  -- 89
        24026 => X"5A",  -- 90
        24027 => X"5A",  -- 90
        24028 => X"55",  -- 85
        24029 => X"4E",  -- 78
        24030 => X"4E",  -- 78
        24031 => X"51",  -- 81
        24032 => X"65",  -- 101
        24033 => X"65",  -- 101
        24034 => X"5A",  -- 90
        24035 => X"45",  -- 69
        24036 => X"3C",  -- 60
        24037 => X"3D",  -- 61
        24038 => X"34",  -- 52
        24039 => X"27",  -- 39
        24040 => X"2A",  -- 42
        24041 => X"2B",  -- 43
        24042 => X"31",  -- 49
        24043 => X"40",  -- 64
        24044 => X"46",  -- 70
        24045 => X"43",  -- 67
        24046 => X"58",  -- 88
        24047 => X"7E",  -- 126
        24048 => X"99",  -- 153
        24049 => X"71",  -- 113
        24050 => X"4D",  -- 77
        24051 => X"41",  -- 65
        24052 => X"3B",  -- 59
        24053 => X"2E",  -- 46
        24054 => X"2F",  -- 47
        24055 => X"41",  -- 65
        24056 => X"51",  -- 81
        24057 => X"4A",  -- 74
        24058 => X"2F",  -- 47
        24059 => X"15",  -- 21
        24060 => X"21",  -- 33
        24061 => X"50",  -- 80
        24062 => X"72",  -- 114
        24063 => X"7A",  -- 122
        24064 => X"73",  -- 115
        24065 => X"87",  -- 135
        24066 => X"93",  -- 147
        24067 => X"9D",  -- 157
        24068 => X"B8",  -- 184
        24069 => X"B8",  -- 184
        24070 => X"C3",  -- 195
        24071 => X"9A",  -- 154
        24072 => X"6C",  -- 108
        24073 => X"3D",  -- 61
        24074 => X"17",  -- 23
        24075 => X"04",  -- 4
        24076 => X"08",  -- 8
        24077 => X"05",  -- 5
        24078 => X"08",  -- 8
        24079 => X"06",  -- 6
        24080 => X"03",  -- 3
        24081 => X"07",  -- 7
        24082 => X"0A",  -- 10
        24083 => X"07",  -- 7
        24084 => X"09",  -- 9
        24085 => X"0D",  -- 13
        24086 => X"14",  -- 20
        24087 => X"17",  -- 23
        24088 => X"2C",  -- 44
        24089 => X"48",  -- 72
        24090 => X"2B",  -- 43
        24091 => X"0A",  -- 10
        24092 => X"06",  -- 6
        24093 => X"2B",  -- 43
        24094 => X"38",  -- 56
        24095 => X"34",  -- 52
        24096 => X"2A",  -- 42
        24097 => X"26",  -- 38
        24098 => X"3A",  -- 58
        24099 => X"13",  -- 19
        24100 => X"15",  -- 21
        24101 => X"09",  -- 9
        24102 => X"22",  -- 34
        24103 => X"3D",  -- 61
        24104 => X"50",  -- 80
        24105 => X"6F",  -- 111
        24106 => X"87",  -- 135
        24107 => X"6D",  -- 109
        24108 => X"2F",  -- 47
        24109 => X"09",  -- 9
        24110 => X"06",  -- 6
        24111 => X"0E",  -- 14
        24112 => X"09",  -- 9
        24113 => X"01",  -- 1
        24114 => X"0D",  -- 13
        24115 => X"0F",  -- 15
        24116 => X"03",  -- 3
        24117 => X"03",  -- 3
        24118 => X"05",  -- 5
        24119 => X"30",  -- 48
        24120 => X"6E",  -- 110
        24121 => X"C0",  -- 192
        24122 => X"C5",  -- 197
        24123 => X"BA",  -- 186
        24124 => X"B8",  -- 184
        24125 => X"A1",  -- 161
        24126 => X"90",  -- 144
        24127 => X"89",  -- 137
        24128 => X"77",  -- 119
        24129 => X"89",  -- 137
        24130 => X"78",  -- 120
        24131 => X"45",  -- 69
        24132 => X"37",  -- 55
        24133 => X"39",  -- 57
        24134 => X"2B",  -- 43
        24135 => X"35",  -- 53
        24136 => X"39",  -- 57
        24137 => X"31",  -- 49
        24138 => X"2A",  -- 42
        24139 => X"2F",  -- 47
        24140 => X"39",  -- 57
        24141 => X"34",  -- 52
        24142 => X"33",  -- 51
        24143 => X"3F",  -- 63
        24144 => X"48",  -- 72
        24145 => X"69",  -- 105
        24146 => X"86",  -- 134
        24147 => X"8E",  -- 142
        24148 => X"8E",  -- 142
        24149 => X"8B",  -- 139
        24150 => X"7F",  -- 127
        24151 => X"6D",  -- 109
        24152 => X"57",  -- 87
        24153 => X"5D",  -- 93
        24154 => X"5C",  -- 92
        24155 => X"50",  -- 80
        24156 => X"49",  -- 73
        24157 => X"52",  -- 82
        24158 => X"61",  -- 97
        24159 => X"6B",  -- 107
        24160 => X"69",  -- 105
        24161 => X"7E",  -- 126
        24162 => X"92",  -- 146
        24163 => X"96",  -- 150
        24164 => X"72",  -- 114
        24165 => X"62",  -- 98
        24166 => X"7D",  -- 125
        24167 => X"80",  -- 128
        24168 => X"7E",  -- 126
        24169 => X"92",  -- 146
        24170 => X"A3",  -- 163
        24171 => X"A3",  -- 163
        24172 => X"9A",  -- 154
        24173 => X"90",  -- 144
        24174 => X"87",  -- 135
        24175 => X"81",  -- 129
        24176 => X"8A",  -- 138
        24177 => X"8A",  -- 138
        24178 => X"82",  -- 130
        24179 => X"71",  -- 113
        24180 => X"63",  -- 99
        24181 => X"5B",  -- 91
        24182 => X"52",  -- 82
        24183 => X"48",  -- 72
        24184 => X"30",  -- 48
        24185 => X"27",  -- 39
        24186 => X"1F",  -- 31
        24187 => X"1F",  -- 31
        24188 => X"20",  -- 32
        24189 => X"28",  -- 40
        24190 => X"47",  -- 71
        24191 => X"69",  -- 105
        24192 => X"7E",  -- 126
        24193 => X"82",  -- 130
        24194 => X"88",  -- 136
        24195 => X"91",  -- 145
        24196 => X"97",  -- 151
        24197 => X"9D",  -- 157
        24198 => X"A9",  -- 169
        24199 => X"B3",  -- 179
        24200 => X"AC",  -- 172
        24201 => X"AD",  -- 173
        24202 => X"AC",  -- 172
        24203 => X"B0",  -- 176
        24204 => X"B3",  -- 179
        24205 => X"B8",  -- 184
        24206 => X"BA",  -- 186
        24207 => X"BB",  -- 187
        24208 => X"BC",  -- 188
        24209 => X"BF",  -- 191
        24210 => X"C3",  -- 195
        24211 => X"C6",  -- 198
        24212 => X"C8",  -- 200
        24213 => X"C9",  -- 201
        24214 => X"CD",  -- 205
        24215 => X"CF",  -- 207
        24216 => X"D1",  -- 209
        24217 => X"CF",  -- 207
        24218 => X"CE",  -- 206
        24219 => X"CB",  -- 203
        24220 => X"C8",  -- 200
        24221 => X"C3",  -- 195
        24222 => X"B8",  -- 184
        24223 => X"AB",  -- 171
        24224 => X"97",  -- 151
        24225 => X"8D",  -- 141
        24226 => X"90",  -- 144
        24227 => X"A1",  -- 161
        24228 => X"B1",  -- 177
        24229 => X"B3",  -- 179
        24230 => X"AF",  -- 175
        24231 => X"AE",  -- 174
        24232 => X"A4",  -- 164
        24233 => X"AF",  -- 175
        24234 => X"B2",  -- 178
        24235 => X"AC",  -- 172
        24236 => X"AC",  -- 172
        24237 => X"B1",  -- 177
        24238 => X"AC",  -- 172
        24239 => X"A0",  -- 160
        24240 => X"97",  -- 151
        24241 => X"9E",  -- 158
        24242 => X"A4",  -- 164
        24243 => X"A4",  -- 164
        24244 => X"9B",  -- 155
        24245 => X"89",  -- 137
        24246 => X"6C",  -- 108
        24247 => X"55",  -- 85
        24248 => X"47",  -- 71
        24249 => X"3E",  -- 62
        24250 => X"40",  -- 64
        24251 => X"54",  -- 84
        24252 => X"70",  -- 112
        24253 => X"84",  -- 132
        24254 => X"91",  -- 145
        24255 => X"97",  -- 151
        24256 => X"9C",  -- 156
        24257 => X"A1",  -- 161
        24258 => X"A6",  -- 166
        24259 => X"A9",  -- 169
        24260 => X"AB",  -- 171
        24261 => X"AE",  -- 174
        24262 => X"B3",  -- 179
        24263 => X"B6",  -- 182
        24264 => X"BC",  -- 188
        24265 => X"C2",  -- 194
        24266 => X"C6",  -- 198
        24267 => X"C8",  -- 200
        24268 => X"C6",  -- 198
        24269 => X"C3",  -- 195
        24270 => X"C1",  -- 193
        24271 => X"C1",  -- 193
        24272 => X"C0",  -- 192
        24273 => X"B0",  -- 176
        24274 => X"71",  -- 113
        24275 => X"29",  -- 41
        24276 => X"24",  -- 36
        24277 => X"50",  -- 80
        24278 => X"75",  -- 117
        24279 => X"7E",  -- 126
        24280 => X"89",  -- 137
        24281 => X"90",  -- 144
        24282 => X"95",  -- 149
        24283 => X"94",  -- 148
        24284 => X"8F",  -- 143
        24285 => X"8D",  -- 141
        24286 => X"93",  -- 147
        24287 => X"99",  -- 153
        24288 => X"95",  -- 149
        24289 => X"A4",  -- 164
        24290 => X"AE",  -- 174
        24291 => X"B2",  -- 178
        24292 => X"B7",  -- 183
        24293 => X"B3",  -- 179
        24294 => X"AE",  -- 174
        24295 => X"AF",  -- 175
        24296 => X"B7",  -- 183
        24297 => X"BB",  -- 187
        24298 => X"BA",  -- 186
        24299 => X"B3",  -- 179
        24300 => X"A7",  -- 167
        24301 => X"A0",  -- 160
        24302 => X"A2",  -- 162
        24303 => X"A6",  -- 166
        24304 => X"AE",  -- 174
        24305 => X"AE",  -- 174
        24306 => X"B1",  -- 177
        24307 => X"B9",  -- 185
        24308 => X"C2",  -- 194
        24309 => X"C3",  -- 195
        24310 => X"B3",  -- 179
        24311 => X"A4",  -- 164
        24312 => X"A3",  -- 163
        24313 => X"A0",  -- 160
        24314 => X"9C",  -- 156
        24315 => X"99",  -- 153
        24316 => X"9E",  -- 158
        24317 => X"A6",  -- 166
        24318 => X"AB",  -- 171
        24319 => X"AB",  -- 171
        24320 => X"98",  -- 152
        24321 => X"9A",  -- 154
        24322 => X"9A",  -- 154
        24323 => X"97",  -- 151
        24324 => X"8C",  -- 140
        24325 => X"7F",  -- 127
        24326 => X"74",  -- 116
        24327 => X"6C",  -- 108
        24328 => X"65",  -- 101
        24329 => X"5E",  -- 94
        24330 => X"5C",  -- 92
        24331 => X"60",  -- 96
        24332 => X"63",  -- 99
        24333 => X"62",  -- 98
        24334 => X"61",  -- 97
        24335 => X"61",  -- 97
        24336 => X"5D",  -- 93
        24337 => X"5C",  -- 92
        24338 => X"58",  -- 88
        24339 => X"57",  -- 87
        24340 => X"59",  -- 89
        24341 => X"58",  -- 88
        24342 => X"56",  -- 86
        24343 => X"54",  -- 84
        24344 => X"52",  -- 82
        24345 => X"50",  -- 80
        24346 => X"52",  -- 82
        24347 => X"54",  -- 84
        24348 => X"52",  -- 82
        24349 => X"4D",  -- 77
        24350 => X"4A",  -- 74
        24351 => X"4A",  -- 74
        24352 => X"53",  -- 83
        24353 => X"5A",  -- 90
        24354 => X"58",  -- 88
        24355 => X"49",  -- 73
        24356 => X"3D",  -- 61
        24357 => X"38",  -- 56
        24358 => X"31",  -- 49
        24359 => X"25",  -- 37
        24360 => X"24",  -- 36
        24361 => X"31",  -- 49
        24362 => X"31",  -- 49
        24363 => X"34",  -- 52
        24364 => X"44",  -- 68
        24365 => X"5E",  -- 94
        24366 => X"7A",  -- 122
        24367 => X"93",  -- 147
        24368 => X"85",  -- 133
        24369 => X"5A",  -- 90
        24370 => X"39",  -- 57
        24371 => X"35",  -- 53
        24372 => X"34",  -- 52
        24373 => X"33",  -- 51
        24374 => X"3D",  -- 61
        24375 => X"4B",  -- 75
        24376 => X"38",  -- 56
        24377 => X"29",  -- 41
        24378 => X"11",  -- 17
        24379 => X"08",  -- 8
        24380 => X"1A",  -- 26
        24381 => X"47",  -- 71
        24382 => X"6E",  -- 110
        24383 => X"80",  -- 128
        24384 => X"7A",  -- 122
        24385 => X"8C",  -- 140
        24386 => X"A3",  -- 163
        24387 => X"AD",  -- 173
        24388 => X"BE",  -- 190
        24389 => X"C1",  -- 193
        24390 => X"B8",  -- 184
        24391 => X"63",  -- 99
        24392 => X"1F",  -- 31
        24393 => X"09",  -- 9
        24394 => X"05",  -- 5
        24395 => X"04",  -- 4
        24396 => X"0E",  -- 14
        24397 => X"04",  -- 4
        24398 => X"06",  -- 6
        24399 => X"04",  -- 4
        24400 => X"01",  -- 1
        24401 => X"05",  -- 5
        24402 => X"07",  -- 7
        24403 => X"07",  -- 7
        24404 => X"0D",  -- 13
        24405 => X"19",  -- 25
        24406 => X"23",  -- 35
        24407 => X"26",  -- 38
        24408 => X"26",  -- 38
        24409 => X"21",  -- 33
        24410 => X"0E",  -- 14
        24411 => X"06",  -- 6
        24412 => X"0B",  -- 11
        24413 => X"3E",  -- 62
        24414 => X"3D",  -- 61
        24415 => X"1F",  -- 31
        24416 => X"28",  -- 40
        24417 => X"1D",  -- 29
        24418 => X"54",  -- 84
        24419 => X"4C",  -- 76
        24420 => X"2E",  -- 46
        24421 => X"15",  -- 21
        24422 => X"3C",  -- 60
        24423 => X"42",  -- 66
        24424 => X"39",  -- 57
        24425 => X"4C",  -- 76
        24426 => X"6C",  -- 108
        24427 => X"78",  -- 120
        24428 => X"5E",  -- 94
        24429 => X"37",  -- 55
        24430 => X"17",  -- 23
        24431 => X"02",  -- 2
        24432 => X"09",  -- 9
        24433 => X"02",  -- 2
        24434 => X"0E",  -- 14
        24435 => X"04",  -- 4
        24436 => X"04",  -- 4
        24437 => X"10",  -- 16
        24438 => X"05",  -- 5
        24439 => X"0C",  -- 12
        24440 => X"2C",  -- 44
        24441 => X"A3",  -- 163
        24442 => X"CB",  -- 203
        24443 => X"BE",  -- 190
        24444 => X"BC",  -- 188
        24445 => X"AD",  -- 173
        24446 => X"A9",  -- 169
        24447 => X"A1",  -- 161
        24448 => X"97",  -- 151
        24449 => X"96",  -- 150
        24450 => X"80",  -- 128
        24451 => X"56",  -- 86
        24452 => X"39",  -- 57
        24453 => X"20",  -- 32
        24454 => X"1C",  -- 28
        24455 => X"46",  -- 70
        24456 => X"6D",  -- 109
        24457 => X"62",  -- 98
        24458 => X"53",  -- 83
        24459 => X"52",  -- 82
        24460 => X"59",  -- 89
        24461 => X"4F",  -- 79
        24462 => X"3E",  -- 62
        24463 => X"38",  -- 56
        24464 => X"44",  -- 68
        24465 => X"50",  -- 80
        24466 => X"62",  -- 98
        24467 => X"73",  -- 115
        24468 => X"84",  -- 132
        24469 => X"91",  -- 145
        24470 => X"98",  -- 152
        24471 => X"9A",  -- 154
        24472 => X"95",  -- 149
        24473 => X"80",  -- 128
        24474 => X"60",  -- 96
        24475 => X"46",  -- 70
        24476 => X"38",  -- 56
        24477 => X"3D",  -- 61
        24478 => X"54",  -- 84
        24479 => X"6C",  -- 108
        24480 => X"6A",  -- 106
        24481 => X"7D",  -- 125
        24482 => X"83",  -- 131
        24483 => X"74",  -- 116
        24484 => X"64",  -- 100
        24485 => X"72",  -- 114
        24486 => X"87",  -- 135
        24487 => X"79",  -- 121
        24488 => X"7D",  -- 125
        24489 => X"8B",  -- 139
        24490 => X"9C",  -- 156
        24491 => X"A1",  -- 161
        24492 => X"9B",  -- 155
        24493 => X"8B",  -- 139
        24494 => X"7B",  -- 123
        24495 => X"70",  -- 112
        24496 => X"79",  -- 121
        24497 => X"84",  -- 132
        24498 => X"86",  -- 134
        24499 => X"7B",  -- 123
        24500 => X"6E",  -- 110
        24501 => X"63",  -- 99
        24502 => X"55",  -- 85
        24503 => X"47",  -- 71
        24504 => X"3B",  -- 59
        24505 => X"26",  -- 38
        24506 => X"1A",  -- 26
        24507 => X"1B",  -- 27
        24508 => X"1D",  -- 29
        24509 => X"25",  -- 37
        24510 => X"46",  -- 70
        24511 => X"6B",  -- 107
        24512 => X"7F",  -- 127
        24513 => X"82",  -- 130
        24514 => X"8D",  -- 141
        24515 => X"9D",  -- 157
        24516 => X"A8",  -- 168
        24517 => X"AB",  -- 171
        24518 => X"AB",  -- 171
        24519 => X"AE",  -- 174
        24520 => X"AF",  -- 175
        24521 => X"AE",  -- 174
        24522 => X"AD",  -- 173
        24523 => X"B0",  -- 176
        24524 => X"B3",  -- 179
        24525 => X"B6",  -- 182
        24526 => X"B9",  -- 185
        24527 => X"BA",  -- 186
        24528 => X"C5",  -- 197
        24529 => X"C7",  -- 199
        24530 => X"C9",  -- 201
        24531 => X"C9",  -- 201
        24532 => X"C7",  -- 199
        24533 => X"C5",  -- 197
        24534 => X"C4",  -- 196
        24535 => X"C4",  -- 196
        24536 => X"C1",  -- 193
        24537 => X"C5",  -- 197
        24538 => X"C6",  -- 198
        24539 => X"C6",  -- 198
        24540 => X"C4",  -- 196
        24541 => X"C2",  -- 194
        24542 => X"BD",  -- 189
        24543 => X"B8",  -- 184
        24544 => X"9F",  -- 159
        24545 => X"97",  -- 151
        24546 => X"98",  -- 152
        24547 => X"A7",  -- 167
        24548 => X"B4",  -- 180
        24549 => X"B6",  -- 182
        24550 => X"B1",  -- 177
        24551 => X"AF",  -- 175
        24552 => X"AF",  -- 175
        24553 => X"B1",  -- 177
        24554 => X"AC",  -- 172
        24555 => X"A7",  -- 167
        24556 => X"AD",  -- 173
        24557 => X"BB",  -- 187
        24558 => X"BC",  -- 188
        24559 => X"B4",  -- 180
        24560 => X"AA",  -- 170
        24561 => X"A6",  -- 166
        24562 => X"A2",  -- 162
        24563 => X"A3",  -- 163
        24564 => X"A4",  -- 164
        24565 => X"95",  -- 149
        24566 => X"6F",  -- 111
        24567 => X"4E",  -- 78
        24568 => X"4B",  -- 75
        24569 => X"44",  -- 68
        24570 => X"44",  -- 68
        24571 => X"50",  -- 80
        24572 => X"67",  -- 103
        24573 => X"7F",  -- 127
        24574 => X"92",  -- 146
        24575 => X"9E",  -- 158
        24576 => X"A3",  -- 163
        24577 => X"A5",  -- 165
        24578 => X"A7",  -- 167
        24579 => X"A8",  -- 168
        24580 => X"A9",  -- 169
        24581 => X"AD",  -- 173
        24582 => X"B3",  -- 179
        24583 => X"B9",  -- 185
        24584 => X"C0",  -- 192
        24585 => X"C4",  -- 196
        24586 => X"C7",  -- 199
        24587 => X"C7",  -- 199
        24588 => X"C6",  -- 198
        24589 => X"C4",  -- 196
        24590 => X"C4",  -- 196
        24591 => X"C4",  -- 196
        24592 => X"B5",  -- 181
        24593 => X"8C",  -- 140
        24594 => X"4A",  -- 74
        24595 => X"22",  -- 34
        24596 => X"36",  -- 54
        24597 => X"62",  -- 98
        24598 => X"78",  -- 120
        24599 => X"79",  -- 121
        24600 => X"86",  -- 134
        24601 => X"91",  -- 145
        24602 => X"9D",  -- 157
        24603 => X"9F",  -- 159
        24604 => X"98",  -- 152
        24605 => X"92",  -- 146
        24606 => X"91",  -- 145
        24607 => X"93",  -- 147
        24608 => X"99",  -- 153
        24609 => X"9D",  -- 157
        24610 => X"A2",  -- 162
        24611 => X"AD",  -- 173
        24612 => X"B3",  -- 179
        24613 => X"AB",  -- 171
        24614 => X"A9",  -- 169
        24615 => X"B3",  -- 179
        24616 => X"AF",  -- 175
        24617 => X"B2",  -- 178
        24618 => X"B0",  -- 176
        24619 => X"AB",  -- 171
        24620 => X"A7",  -- 167
        24621 => X"A5",  -- 165
        24622 => X"A8",  -- 168
        24623 => X"AB",  -- 171
        24624 => X"AE",  -- 174
        24625 => X"B0",  -- 176
        24626 => X"B4",  -- 180
        24627 => X"BA",  -- 186
        24628 => X"C3",  -- 195
        24629 => X"C5",  -- 197
        24630 => X"BA",  -- 186
        24631 => X"AE",  -- 174
        24632 => X"A1",  -- 161
        24633 => X"9F",  -- 159
        24634 => X"9D",  -- 157
        24635 => X"9E",  -- 158
        24636 => X"9F",  -- 159
        24637 => X"A1",  -- 161
        24638 => X"A5",  -- 165
        24639 => X"A8",  -- 168
        24640 => X"88",  -- 136
        24641 => X"89",  -- 137
        24642 => X"8A",  -- 138
        24643 => X"86",  -- 134
        24644 => X"7F",  -- 127
        24645 => X"74",  -- 116
        24646 => X"6A",  -- 106
        24647 => X"65",  -- 101
        24648 => X"5D",  -- 93
        24649 => X"53",  -- 83
        24650 => X"4C",  -- 76
        24651 => X"4F",  -- 79
        24652 => X"54",  -- 84
        24653 => X"55",  -- 85
        24654 => X"57",  -- 87
        24655 => X"58",  -- 88
        24656 => X"55",  -- 85
        24657 => X"53",  -- 83
        24658 => X"53",  -- 83
        24659 => X"52",  -- 82
        24660 => X"53",  -- 83
        24661 => X"54",  -- 84
        24662 => X"52",  -- 82
        24663 => X"50",  -- 80
        24664 => X"4F",  -- 79
        24665 => X"4B",  -- 75
        24666 => X"49",  -- 73
        24667 => X"4D",  -- 77
        24668 => X"4F",  -- 79
        24669 => X"4C",  -- 76
        24670 => X"47",  -- 71
        24671 => X"44",  -- 68
        24672 => X"44",  -- 68
        24673 => X"4E",  -- 78
        24674 => X"53",  -- 83
        24675 => X"4B",  -- 75
        24676 => X"3E",  -- 62
        24677 => X"33",  -- 51
        24678 => X"2C",  -- 44
        24679 => X"27",  -- 39
        24680 => X"28",  -- 40
        24681 => X"3F",  -- 63
        24682 => X"4F",  -- 79
        24683 => X"5C",  -- 92
        24684 => X"7C",  -- 124
        24685 => X"99",  -- 153
        24686 => X"9D",  -- 157
        24687 => X"97",  -- 151
        24688 => X"53",  -- 83
        24689 => X"3B",  -- 59
        24690 => X"2B",  -- 43
        24691 => X"2A",  -- 42
        24692 => X"38",  -- 56
        24693 => X"51",  -- 81
        24694 => X"57",  -- 87
        24695 => X"49",  -- 73
        24696 => X"21",  -- 33
        24697 => X"10",  -- 16
        24698 => X"07",  -- 7
        24699 => X"15",  -- 21
        24700 => X"37",  -- 55
        24701 => X"5C",  -- 92
        24702 => X"76",  -- 118
        24703 => X"84",  -- 132
        24704 => X"97",  -- 151
        24705 => X"9E",  -- 158
        24706 => X"AD",  -- 173
        24707 => X"BA",  -- 186
        24708 => X"C8",  -- 200
        24709 => X"C1",  -- 193
        24710 => X"88",  -- 136
        24711 => X"1E",  -- 30
        24712 => X"05",  -- 5
        24713 => X"01",  -- 1
        24714 => X"02",  -- 2
        24715 => X"04",  -- 4
        24716 => X"07",  -- 7
        24717 => X"01",  -- 1
        24718 => X"02",  -- 2
        24719 => X"07",  -- 7
        24720 => X"02",  -- 2
        24721 => X"04",  -- 4
        24722 => X"0C",  -- 12
        24723 => X"1C",  -- 28
        24724 => X"2D",  -- 45
        24725 => X"38",  -- 56
        24726 => X"36",  -- 54
        24727 => X"2F",  -- 47
        24728 => X"21",  -- 33
        24729 => X"12",  -- 18
        24730 => X"0B",  -- 11
        24731 => X"14",  -- 20
        24732 => X"27",  -- 39
        24733 => X"58",  -- 88
        24734 => X"41",  -- 65
        24735 => X"18",  -- 24
        24736 => X"41",  -- 65
        24737 => X"19",  -- 25
        24738 => X"2C",  -- 44
        24739 => X"4A",  -- 74
        24740 => X"59",  -- 89
        24741 => X"40",  -- 64
        24742 => X"5C",  -- 92
        24743 => X"7C",  -- 124
        24744 => X"57",  -- 87
        24745 => X"56",  -- 86
        24746 => X"68",  -- 104
        24747 => X"80",  -- 128
        24748 => X"84",  -- 132
        24749 => X"6B",  -- 107
        24750 => X"3F",  -- 63
        24751 => X"17",  -- 23
        24752 => X"11",  -- 17
        24753 => X"02",  -- 2
        24754 => X"00",  -- 0
        24755 => X"03",  -- 3
        24756 => X"0C",  -- 12
        24757 => X"0F",  -- 15
        24758 => X"01",  -- 1
        24759 => X"01",  -- 1
        24760 => X"10",  -- 16
        24761 => X"7F",  -- 127
        24762 => X"C4",  -- 196
        24763 => X"C0",  -- 192
        24764 => X"C4",  -- 196
        24765 => X"C0",  -- 192
        24766 => X"BD",  -- 189
        24767 => X"AB",  -- 171
        24768 => X"A0",  -- 160
        24769 => X"96",  -- 150
        24770 => X"93",  -- 147
        24771 => X"62",  -- 98
        24772 => X"20",  -- 32
        24773 => X"15",  -- 21
        24774 => X"22",  -- 34
        24775 => X"2C",  -- 44
        24776 => X"64",  -- 100
        24777 => X"71",  -- 113
        24778 => X"72",  -- 114
        24779 => X"6A",  -- 106
        24780 => X"61",  -- 97
        24781 => X"4E",  -- 78
        24782 => X"32",  -- 50
        24783 => X"25",  -- 37
        24784 => X"31",  -- 49
        24785 => X"37",  -- 55
        24786 => X"4C",  -- 76
        24787 => X"6E",  -- 110
        24788 => X"87",  -- 135
        24789 => X"8C",  -- 140
        24790 => X"8A",  -- 138
        24791 => X"87",  -- 135
        24792 => X"8E",  -- 142
        24793 => X"82",  -- 130
        24794 => X"7B",  -- 123
        24795 => X"76",  -- 118
        24796 => X"6A",  -- 106
        24797 => X"5A",  -- 90
        24798 => X"57",  -- 87
        24799 => X"5D",  -- 93
        24800 => X"63",  -- 99
        24801 => X"82",  -- 130
        24802 => X"85",  -- 133
        24803 => X"6D",  -- 109
        24804 => X"6B",  -- 107
        24805 => X"80",  -- 128
        24806 => X"83",  -- 131
        24807 => X"73",  -- 115
        24808 => X"6E",  -- 110
        24809 => X"80",  -- 128
        24810 => X"97",  -- 151
        24811 => X"A3",  -- 163
        24812 => X"9D",  -- 157
        24813 => X"8C",  -- 140
        24814 => X"80",  -- 128
        24815 => X"7B",  -- 123
        24816 => X"79",  -- 121
        24817 => X"84",  -- 132
        24818 => X"88",  -- 136
        24819 => X"7B",  -- 123
        24820 => X"6E",  -- 110
        24821 => X"61",  -- 97
        24822 => X"52",  -- 82
        24823 => X"41",  -- 65
        24824 => X"49",  -- 73
        24825 => X"30",  -- 48
        24826 => X"1F",  -- 31
        24827 => X"1D",  -- 29
        24828 => X"1C",  -- 28
        24829 => X"22",  -- 34
        24830 => X"3F",  -- 63
        24831 => X"64",  -- 100
        24832 => X"8C",  -- 140
        24833 => X"8D",  -- 141
        24834 => X"95",  -- 149
        24835 => X"A0",  -- 160
        24836 => X"AA",  -- 170
        24837 => X"AD",  -- 173
        24838 => X"AF",  -- 175
        24839 => X"AE",  -- 174
        24840 => X"B7",  -- 183
        24841 => X"B8",  -- 184
        24842 => X"B7",  -- 183
        24843 => X"B7",  -- 183
        24844 => X"B9",  -- 185
        24845 => X"BC",  -- 188
        24846 => X"BD",  -- 189
        24847 => X"BE",  -- 190
        24848 => X"C3",  -- 195
        24849 => X"C5",  -- 197
        24850 => X"C7",  -- 199
        24851 => X"C7",  -- 199
        24852 => X"C7",  -- 199
        24853 => X"C4",  -- 196
        24854 => X"C3",  -- 195
        24855 => X"C1",  -- 193
        24856 => X"C1",  -- 193
        24857 => X"C7",  -- 199
        24858 => X"CC",  -- 204
        24859 => X"CC",  -- 204
        24860 => X"CB",  -- 203
        24861 => X"CA",  -- 202
        24862 => X"C8",  -- 200
        24863 => X"C2",  -- 194
        24864 => X"AA",  -- 170
        24865 => X"A1",  -- 161
        24866 => X"A0",  -- 160
        24867 => X"A8",  -- 168
        24868 => X"B3",  -- 179
        24869 => X"B6",  -- 182
        24870 => X"B4",  -- 180
        24871 => X"B1",  -- 177
        24872 => X"AF",  -- 175
        24873 => X"AE",  -- 174
        24874 => X"AA",  -- 170
        24875 => X"A9",  -- 169
        24876 => X"AF",  -- 175
        24877 => X"B7",  -- 183
        24878 => X"B2",  -- 178
        24879 => X"AA",  -- 170
        24880 => X"99",  -- 153
        24881 => X"96",  -- 150
        24882 => X"94",  -- 148
        24883 => X"96",  -- 150
        24884 => X"98",  -- 152
        24885 => X"91",  -- 145
        24886 => X"7A",  -- 122
        24887 => X"66",  -- 102
        24888 => X"59",  -- 89
        24889 => X"54",  -- 84
        24890 => X"51",  -- 81
        24891 => X"5A",  -- 90
        24892 => X"6F",  -- 111
        24893 => X"87",  -- 135
        24894 => X"9B",  -- 155
        24895 => X"A5",  -- 165
        24896 => X"A5",  -- 165
        24897 => X"A5",  -- 165
        24898 => X"A6",  -- 166
        24899 => X"A6",  -- 166
        24900 => X"A9",  -- 169
        24901 => X"AF",  -- 175
        24902 => X"B8",  -- 184
        24903 => X"BD",  -- 189
        24904 => X"BC",  -- 188
        24905 => X"C1",  -- 193
        24906 => X"C5",  -- 197
        24907 => X"C4",  -- 196
        24908 => X"C5",  -- 197
        24909 => X"C6",  -- 198
        24910 => X"C8",  -- 200
        24911 => X"C7",  -- 199
        24912 => X"B5",  -- 181
        24913 => X"67",  -- 103
        24914 => X"28",  -- 40
        24915 => X"2B",  -- 43
        24916 => X"4C",  -- 76
        24917 => X"66",  -- 102
        24918 => X"78",  -- 120
        24919 => X"86",  -- 134
        24920 => X"9D",  -- 157
        24921 => X"A2",  -- 162
        24922 => X"A4",  -- 164
        24923 => X"A0",  -- 160
        24924 => X"9C",  -- 156
        24925 => X"9A",  -- 154
        24926 => X"9D",  -- 157
        24927 => X"A2",  -- 162
        24928 => X"A7",  -- 167
        24929 => X"A4",  -- 164
        24930 => X"A1",  -- 161
        24931 => X"A8",  -- 168
        24932 => X"AE",  -- 174
        24933 => X"A7",  -- 167
        24934 => X"A8",  -- 168
        24935 => X"BA",  -- 186
        24936 => X"B4",  -- 180
        24937 => X"B1",  -- 177
        24938 => X"A8",  -- 168
        24939 => X"9E",  -- 158
        24940 => X"9B",  -- 155
        24941 => X"9F",  -- 159
        24942 => X"A6",  -- 166
        24943 => X"AA",  -- 170
        24944 => X"AC",  -- 172
        24945 => X"B0",  -- 176
        24946 => X"B7",  -- 183
        24947 => X"BE",  -- 190
        24948 => X"C4",  -- 196
        24949 => X"C6",  -- 198
        24950 => X"BE",  -- 190
        24951 => X"B4",  -- 180
        24952 => X"A4",  -- 164
        24953 => X"A1",  -- 161
        24954 => X"A1",  -- 161
        24955 => X"A3",  -- 163
        24956 => X"A3",  -- 163
        24957 => X"A0",  -- 160
        24958 => X"A3",  -- 163
        24959 => X"A8",  -- 168
        24960 => X"79",  -- 121
        24961 => X"7A",  -- 122
        24962 => X"79",  -- 121
        24963 => X"76",  -- 118
        24964 => X"70",  -- 112
        24965 => X"6C",  -- 108
        24966 => X"69",  -- 105
        24967 => X"69",  -- 105
        24968 => X"63",  -- 99
        24969 => X"58",  -- 88
        24970 => X"4F",  -- 79
        24971 => X"4F",  -- 79
        24972 => X"53",  -- 83
        24973 => X"56",  -- 86
        24974 => X"57",  -- 87
        24975 => X"57",  -- 87
        24976 => X"59",  -- 89
        24977 => X"59",  -- 89
        24978 => X"5A",  -- 90
        24979 => X"59",  -- 89
        24980 => X"59",  -- 89
        24981 => X"59",  -- 89
        24982 => X"59",  -- 89
        24983 => X"59",  -- 89
        24984 => X"57",  -- 87
        24985 => X"51",  -- 81
        24986 => X"4D",  -- 77
        24987 => X"4F",  -- 79
        24988 => X"50",  -- 80
        24989 => X"4C",  -- 76
        24990 => X"49",  -- 73
        24991 => X"48",  -- 72
        24992 => X"43",  -- 67
        24993 => X"43",  -- 67
        24994 => X"44",  -- 68
        24995 => X"42",  -- 66
        24996 => X"37",  -- 55
        24997 => X"2E",  -- 46
        24998 => X"30",  -- 48
        24999 => X"37",  -- 55
        25000 => X"4C",  -- 76
        25001 => X"51",  -- 81
        25002 => X"5B",  -- 91
        25003 => X"77",  -- 119
        25004 => X"9D",  -- 157
        25005 => X"9E",  -- 158
        25006 => X"71",  -- 113
        25007 => X"48",  -- 72
        25008 => X"3A",  -- 58
        25009 => X"26",  -- 38
        25010 => X"20",  -- 32
        25011 => X"2C",  -- 44
        25012 => X"47",  -- 71
        25013 => X"65",  -- 101
        25014 => X"5D",  -- 93
        25015 => X"35",  -- 53
        25016 => X"17",  -- 23
        25017 => X"06",  -- 6
        25018 => X"07",  -- 7
        25019 => X"2A",  -- 42
        25020 => X"5C",  -- 92
        25021 => X"7E",  -- 126
        25022 => X"8B",  -- 139
        25023 => X"8F",  -- 143
        25024 => X"AF",  -- 175
        25025 => X"B8",  -- 184
        25026 => X"BA",  -- 186
        25027 => X"C5",  -- 197
        25028 => X"D4",  -- 212
        25029 => X"B6",  -- 182
        25030 => X"4D",  -- 77
        25031 => X"02",  -- 2
        25032 => X"0A",  -- 10
        25033 => X"09",  -- 9
        25034 => X"05",  -- 5
        25035 => X"08",  -- 8
        25036 => X"02",  -- 2
        25037 => X"04",  -- 4
        25038 => X"07",  -- 7
        25039 => X"11",  -- 17
        25040 => X"19",  -- 25
        25041 => X"27",  -- 39
        25042 => X"42",  -- 66
        25043 => X"5D",  -- 93
        25044 => X"69",  -- 105
        25045 => X"5F",  -- 95
        25046 => X"4C",  -- 76
        25047 => X"3D",  -- 61
        25048 => X"3E",  -- 62
        25049 => X"3A",  -- 58
        25050 => X"33",  -- 51
        25051 => X"3C",  -- 60
        25052 => X"54",  -- 84
        25053 => X"69",  -- 105
        25054 => X"37",  -- 55
        25055 => X"1B",  -- 27
        25056 => X"54",  -- 84
        25057 => X"35",  -- 53
        25058 => X"14",  -- 20
        25059 => X"1D",  -- 29
        25060 => X"4F",  -- 79
        25061 => X"54",  -- 84
        25062 => X"66",  -- 102
        25063 => X"8B",  -- 139
        25064 => X"74",  -- 116
        25065 => X"79",  -- 121
        25066 => X"86",  -- 134
        25067 => X"8D",  -- 141
        25068 => X"8C",  -- 140
        25069 => X"87",  -- 135
        25070 => X"74",  -- 116
        25071 => X"5A",  -- 90
        25072 => X"3C",  -- 60
        25073 => X"1F",  -- 31
        25074 => X"04",  -- 4
        25075 => X"07",  -- 7
        25076 => X"09",  -- 9
        25077 => X"01",  -- 1
        25078 => X"07",  -- 7
        25079 => X"0E",  -- 14
        25080 => X"11",  -- 17
        25081 => X"61",  -- 97
        25082 => X"BF",  -- 191
        25083 => X"CA",  -- 202
        25084 => X"CC",  -- 204
        25085 => X"C9",  -- 201
        25086 => X"C5",  -- 197
        25087 => X"B4",  -- 180
        25088 => X"AE",  -- 174
        25089 => X"98",  -- 152
        25090 => X"93",  -- 147
        25091 => X"76",  -- 118
        25092 => X"53",  -- 83
        25093 => X"4D",  -- 77
        25094 => X"39",  -- 57
        25095 => X"1C",  -- 28
        25096 => X"2A",  -- 42
        25097 => X"56",  -- 86
        25098 => X"73",  -- 115
        25099 => X"70",  -- 112
        25100 => X"69",  -- 105
        25101 => X"5A",  -- 90
        25102 => X"45",  -- 69
        25103 => X"39",  -- 57
        25104 => X"35",  -- 53
        25105 => X"34",  -- 52
        25106 => X"41",  -- 65
        25107 => X"64",  -- 100
        25108 => X"88",  -- 136
        25109 => X"9C",  -- 156
        25110 => X"A2",  -- 162
        25111 => X"A2",  -- 162
        25112 => X"97",  -- 151
        25113 => X"8A",  -- 138
        25114 => X"74",  -- 116
        25115 => X"5F",  -- 95
        25116 => X"4D",  -- 77
        25117 => X"44",  -- 68
        25118 => X"45",  -- 69
        25119 => X"4B",  -- 75
        25120 => X"58",  -- 88
        25121 => X"75",  -- 117
        25122 => X"74",  -- 116
        25123 => X"62",  -- 98
        25124 => X"77",  -- 119
        25125 => X"8C",  -- 140
        25126 => X"81",  -- 129
        25127 => X"78",  -- 120
        25128 => X"67",  -- 103
        25129 => X"74",  -- 116
        25130 => X"8B",  -- 139
        25131 => X"9D",  -- 157
        25132 => X"9C",  -- 156
        25133 => X"8F",  -- 143
        25134 => X"85",  -- 133
        25135 => X"81",  -- 129
        25136 => X"87",  -- 135
        25137 => X"90",  -- 144
        25138 => X"8E",  -- 142
        25139 => X"7F",  -- 127
        25140 => X"71",  -- 113
        25141 => X"6A",  -- 106
        25142 => X"5D",  -- 93
        25143 => X"4E",  -- 78
        25144 => X"45",  -- 69
        25145 => X"32",  -- 50
        25146 => X"24",  -- 36
        25147 => X"1D",  -- 29
        25148 => X"16",  -- 22
        25149 => X"15",  -- 21
        25150 => X"2D",  -- 45
        25151 => X"4F",  -- 79
        25152 => X"8D",  -- 141
        25153 => X"91",  -- 145
        25154 => X"96",  -- 150
        25155 => X"99",  -- 153
        25156 => X"9E",  -- 158
        25157 => X"A7",  -- 167
        25158 => X"AF",  -- 175
        25159 => X"B3",  -- 179
        25160 => X"BA",  -- 186
        25161 => X"BB",  -- 187
        25162 => X"BD",  -- 189
        25163 => X"BC",  -- 188
        25164 => X"BA",  -- 186
        25165 => X"BC",  -- 188
        25166 => X"BE",  -- 190
        25167 => X"C2",  -- 194
        25168 => X"C0",  -- 192
        25169 => X"C0",  -- 192
        25170 => X"C0",  -- 192
        25171 => X"C2",  -- 194
        25172 => X"C3",  -- 195
        25173 => X"C3",  -- 195
        25174 => X"C2",  -- 194
        25175 => X"C2",  -- 194
        25176 => X"C6",  -- 198
        25177 => X"CA",  -- 202
        25178 => X"CF",  -- 207
        25179 => X"D1",  -- 209
        25180 => X"D2",  -- 210
        25181 => X"CE",  -- 206
        25182 => X"C5",  -- 197
        25183 => X"BB",  -- 187
        25184 => X"A9",  -- 169
        25185 => X"9E",  -- 158
        25186 => X"98",  -- 152
        25187 => X"9F",  -- 159
        25188 => X"AA",  -- 170
        25189 => X"B3",  -- 179
        25190 => X"B6",  -- 182
        25191 => X"B8",  -- 184
        25192 => X"B0",  -- 176
        25193 => X"AF",  -- 175
        25194 => X"B0",  -- 176
        25195 => X"B1",  -- 177
        25196 => X"B2",  -- 178
        25197 => X"AC",  -- 172
        25198 => X"A4",  -- 164
        25199 => X"9B",  -- 155
        25200 => X"97",  -- 151
        25201 => X"9A",  -- 154
        25202 => X"99",  -- 153
        25203 => X"91",  -- 145
        25204 => X"87",  -- 135
        25205 => X"7B",  -- 123
        25206 => X"6A",  -- 106
        25207 => X"5F",  -- 95
        25208 => X"49",  -- 73
        25209 => X"44",  -- 68
        25210 => X"45",  -- 69
        25211 => X"55",  -- 85
        25212 => X"70",  -- 112
        25213 => X"8A",  -- 138
        25214 => X"99",  -- 153
        25215 => X"9C",  -- 156
        25216 => X"9E",  -- 158
        25217 => X"A2",  -- 162
        25218 => X"A4",  -- 164
        25219 => X"A8",  -- 168
        25220 => X"AC",  -- 172
        25221 => X"B2",  -- 178
        25222 => X"BC",  -- 188
        25223 => X"C3",  -- 195
        25224 => X"C2",  -- 194
        25225 => X"C5",  -- 197
        25226 => X"C5",  -- 197
        25227 => X"C3",  -- 195
        25228 => X"C4",  -- 196
        25229 => X"C5",  -- 197
        25230 => X"C1",  -- 193
        25231 => X"BA",  -- 186
        25232 => X"9F",  -- 159
        25233 => X"4B",  -- 75
        25234 => X"1D",  -- 29
        25235 => X"35",  -- 53
        25236 => X"56",  -- 86
        25237 => X"6E",  -- 110
        25238 => X"83",  -- 131
        25239 => X"8F",  -- 143
        25240 => X"A2",  -- 162
        25241 => X"9E",  -- 158
        25242 => X"97",  -- 151
        25243 => X"92",  -- 146
        25244 => X"8F",  -- 143
        25245 => X"91",  -- 145
        25246 => X"96",  -- 150
        25247 => X"9A",  -- 154
        25248 => X"9C",  -- 156
        25249 => X"9E",  -- 158
        25250 => X"9B",  -- 155
        25251 => X"9F",  -- 159
        25252 => X"A6",  -- 166
        25253 => X"A5",  -- 165
        25254 => X"A4",  -- 164
        25255 => X"AE",  -- 174
        25256 => X"BA",  -- 186
        25257 => X"B8",  -- 184
        25258 => X"AF",  -- 175
        25259 => X"A1",  -- 161
        25260 => X"98",  -- 152
        25261 => X"9B",  -- 155
        25262 => X"A2",  -- 162
        25263 => X"A6",  -- 166
        25264 => X"A9",  -- 169
        25265 => X"B2",  -- 178
        25266 => X"BA",  -- 186
        25267 => X"C2",  -- 194
        25268 => X"C8",  -- 200
        25269 => X"C8",  -- 200
        25270 => X"C1",  -- 193
        25271 => X"B9",  -- 185
        25272 => X"AA",  -- 170
        25273 => X"A3",  -- 163
        25274 => X"A0",  -- 160
        25275 => X"A4",  -- 164
        25276 => X"A5",  -- 165
        25277 => X"A1",  -- 161
        25278 => X"A2",  -- 162
        25279 => X"A8",  -- 168
        25280 => X"70",  -- 112
        25281 => X"70",  -- 112
        25282 => X"6C",  -- 108
        25283 => X"69",  -- 105
        25284 => X"66",  -- 102
        25285 => X"67",  -- 103
        25286 => X"6B",  -- 107
        25287 => X"6D",  -- 109
        25288 => X"6C",  -- 108
        25289 => X"60",  -- 96
        25290 => X"55",  -- 85
        25291 => X"57",  -- 87
        25292 => X"5A",  -- 90
        25293 => X"5D",  -- 93
        25294 => X"5D",  -- 93
        25295 => X"5F",  -- 95
        25296 => X"60",  -- 96
        25297 => X"61",  -- 97
        25298 => X"62",  -- 98
        25299 => X"62",  -- 98
        25300 => X"63",  -- 99
        25301 => X"63",  -- 99
        25302 => X"62",  -- 98
        25303 => X"61",  -- 97
        25304 => X"5C",  -- 92
        25305 => X"57",  -- 87
        25306 => X"55",  -- 85
        25307 => X"57",  -- 87
        25308 => X"57",  -- 87
        25309 => X"54",  -- 84
        25310 => X"54",  -- 84
        25311 => X"56",  -- 86
        25312 => X"4A",  -- 74
        25313 => X"40",  -- 64
        25314 => X"37",  -- 55
        25315 => X"34",  -- 52
        25316 => X"2E",  -- 46
        25317 => X"2D",  -- 45
        25318 => X"3A",  -- 58
        25319 => X"4C",  -- 76
        25320 => X"52",  -- 82
        25321 => X"68",  -- 104
        25322 => X"84",  -- 132
        25323 => X"9B",  -- 155
        25324 => X"9B",  -- 155
        25325 => X"77",  -- 119
        25326 => X"51",  -- 81
        25327 => X"45",  -- 69
        25328 => X"36",  -- 54
        25329 => X"26",  -- 38
        25330 => X"31",  -- 49
        25331 => X"4D",  -- 77
        25332 => X"5C",  -- 92
        25333 => X"5E",  -- 94
        25334 => X"46",  -- 70
        25335 => X"20",  -- 32
        25336 => X"0C",  -- 12
        25337 => X"06",  -- 6
        25338 => X"10",  -- 16
        25339 => X"38",  -- 56
        25340 => X"6A",  -- 106
        25341 => X"8C",  -- 140
        25342 => X"9C",  -- 156
        25343 => X"A2",  -- 162
        25344 => X"AD",  -- 173
        25345 => X"C3",  -- 195
        25346 => X"C1",  -- 193
        25347 => X"CC",  -- 204
        25348 => X"DF",  -- 223
        25349 => X"AF",  -- 175
        25350 => X"2C",  -- 44
        25351 => X"0F",  -- 15
        25352 => X"02",  -- 2
        25353 => X"07",  -- 7
        25354 => X"07",  -- 7
        25355 => X"1A",  -- 26
        25356 => X"1F",  -- 31
        25357 => X"37",  -- 55
        25358 => X"3E",  -- 62
        25359 => X"4C",  -- 76
        25360 => X"6A",  -- 106
        25361 => X"6B",  -- 107
        25362 => X"70",  -- 112
        25363 => X"72",  -- 114
        25364 => X"6B",  -- 107
        25365 => X"67",  -- 103
        25366 => X"71",  -- 113
        25367 => X"7E",  -- 126
        25368 => X"73",  -- 115
        25369 => X"7B",  -- 123
        25370 => X"6A",  -- 106
        25371 => X"62",  -- 98
        25372 => X"70",  -- 112
        25373 => X"69",  -- 105
        25374 => X"22",  -- 34
        25375 => X"1C",  -- 28
        25376 => X"58",  -- 88
        25377 => X"51",  -- 81
        25378 => X"31",  -- 49
        25379 => X"12",  -- 18
        25380 => X"0F",  -- 15
        25381 => X"43",  -- 67
        25382 => X"74",  -- 116
        25383 => X"6C",  -- 108
        25384 => X"71",  -- 113
        25385 => X"85",  -- 133
        25386 => X"93",  -- 147
        25387 => X"8B",  -- 139
        25388 => X"83",  -- 131
        25389 => X"90",  -- 144
        25390 => X"98",  -- 152
        25391 => X"8D",  -- 141
        25392 => X"87",  -- 135
        25393 => X"85",  -- 133
        25394 => X"5B",  -- 91
        25395 => X"3C",  -- 60
        25396 => X"26",  -- 38
        25397 => X"17",  -- 23
        25398 => X"18",  -- 24
        25399 => X"03",  -- 3
        25400 => X"14",  -- 20
        25401 => X"4C",  -- 76
        25402 => X"BF",  -- 191
        25403 => X"D6",  -- 214
        25404 => X"D1",  -- 209
        25405 => X"CD",  -- 205
        25406 => X"CE",  -- 206
        25407 => X"C5",  -- 197
        25408 => X"AD",  -- 173
        25409 => X"A3",  -- 163
        25410 => X"A5",  -- 165
        25411 => X"AA",  -- 170
        25412 => X"8C",  -- 140
        25413 => X"35",  -- 53
        25414 => X"05",  -- 5
        25415 => X"0D",  -- 13
        25416 => X"21",  -- 33
        25417 => X"58",  -- 88
        25418 => X"7E",  -- 126
        25419 => X"80",  -- 128
        25420 => X"7A",  -- 122
        25421 => X"71",  -- 113
        25422 => X"60",  -- 96
        25423 => X"50",  -- 80
        25424 => X"2D",  -- 45
        25425 => X"28",  -- 40
        25426 => X"2C",  -- 44
        25427 => X"47",  -- 71
        25428 => X"6E",  -- 110
        25429 => X"90",  -- 144
        25430 => X"A3",  -- 163
        25431 => X"A6",  -- 166
        25432 => X"A9",  -- 169
        25433 => X"AD",  -- 173
        25434 => X"A4",  -- 164
        25435 => X"8B",  -- 139
        25436 => X"6E",  -- 110
        25437 => X"5A",  -- 90
        25438 => X"46",  -- 70
        25439 => X"37",  -- 55
        25440 => X"5A",  -- 90
        25441 => X"5F",  -- 95
        25442 => X"4A",  -- 74
        25443 => X"48",  -- 72
        25444 => X"81",  -- 129
        25445 => X"9F",  -- 159
        25446 => X"85",  -- 133
        25447 => X"7B",  -- 123
        25448 => X"6F",  -- 111
        25449 => X"73",  -- 115
        25450 => X"81",  -- 129
        25451 => X"94",  -- 148
        25452 => X"98",  -- 152
        25453 => X"8A",  -- 138
        25454 => X"78",  -- 120
        25455 => X"6D",  -- 109
        25456 => X"81",  -- 129
        25457 => X"8E",  -- 142
        25458 => X"93",  -- 147
        25459 => X"8A",  -- 138
        25460 => X"82",  -- 130
        25461 => X"7E",  -- 126
        25462 => X"6F",  -- 111
        25463 => X"5E",  -- 94
        25464 => X"4A",  -- 74
        25465 => X"3D",  -- 61
        25466 => X"33",  -- 51
        25467 => X"2C",  -- 44
        25468 => X"1C",  -- 28
        25469 => X"16",  -- 22
        25470 => X"2D",  -- 45
        25471 => X"4B",  -- 75
        25472 => X"70",  -- 112
        25473 => X"82",  -- 130
        25474 => X"94",  -- 148
        25475 => X"9C",  -- 156
        25476 => X"A0",  -- 160
        25477 => X"A8",  -- 168
        25478 => X"B0",  -- 176
        25479 => X"B2",  -- 178
        25480 => X"B4",  -- 180
        25481 => X"B8",  -- 184
        25482 => X"BA",  -- 186
        25483 => X"B8",  -- 184
        25484 => X"B7",  -- 183
        25485 => X"B7",  -- 183
        25486 => X"BB",  -- 187
        25487 => X"BF",  -- 191
        25488 => X"C3",  -- 195
        25489 => X"C1",  -- 193
        25490 => X"BE",  -- 190
        25491 => X"BC",  -- 188
        25492 => X"BD",  -- 189
        25493 => X"BD",  -- 189
        25494 => X"BD",  -- 189
        25495 => X"BC",  -- 188
        25496 => X"BA",  -- 186
        25497 => X"C0",  -- 192
        25498 => X"C6",  -- 198
        25499 => X"CB",  -- 203
        25500 => X"D0",  -- 208
        25501 => X"CC",  -- 204
        25502 => X"BD",  -- 189
        25503 => X"AE",  -- 174
        25504 => X"9B",  -- 155
        25505 => X"91",  -- 145
        25506 => X"8A",  -- 138
        25507 => X"90",  -- 144
        25508 => X"9D",  -- 157
        25509 => X"AB",  -- 171
        25510 => X"B5",  -- 181
        25511 => X"B9",  -- 185
        25512 => X"B9",  -- 185
        25513 => X"B6",  -- 182
        25514 => X"B4",  -- 180
        25515 => X"B3",  -- 179
        25516 => X"B0",  -- 176
        25517 => X"AB",  -- 171
        25518 => X"AB",  -- 171
        25519 => X"AD",  -- 173
        25520 => X"A7",  -- 167
        25521 => X"A0",  -- 160
        25522 => X"97",  -- 151
        25523 => X"94",  -- 148
        25524 => X"91",  -- 145
        25525 => X"85",  -- 133
        25526 => X"6C",  -- 108
        25527 => X"53",  -- 83
        25528 => X"37",  -- 55
        25529 => X"34",  -- 52
        25530 => X"39",  -- 57
        25531 => X"52",  -- 82
        25532 => X"75",  -- 117
        25533 => X"93",  -- 147
        25534 => X"9D",  -- 157
        25535 => X"9A",  -- 154
        25536 => X"98",  -- 152
        25537 => X"9C",  -- 156
        25538 => X"A3",  -- 163
        25539 => X"A8",  -- 168
        25540 => X"AF",  -- 175
        25541 => X"B7",  -- 183
        25542 => X"C1",  -- 193
        25543 => X"C8",  -- 200
        25544 => X"CC",  -- 204
        25545 => X"CD",  -- 205
        25546 => X"CB",  -- 203
        25547 => X"C7",  -- 199
        25548 => X"C2",  -- 194
        25549 => X"BE",  -- 190
        25550 => X"B4",  -- 180
        25551 => X"AA",  -- 170
        25552 => X"6B",  -- 107
        25553 => X"31",  -- 49
        25554 => X"20",  -- 32
        25555 => X"3F",  -- 63
        25556 => X"5F",  -- 95
        25557 => X"81",  -- 129
        25558 => X"92",  -- 146
        25559 => X"89",  -- 137
        25560 => X"96",  -- 150
        25561 => X"98",  -- 152
        25562 => X"9A",  -- 154
        25563 => X"9C",  -- 156
        25564 => X"9C",  -- 156
        25565 => X"96",  -- 150
        25566 => X"8E",  -- 142
        25567 => X"87",  -- 135
        25568 => X"8C",  -- 140
        25569 => X"9A",  -- 154
        25570 => X"A0",  -- 160
        25571 => X"A5",  -- 165
        25572 => X"AD",  -- 173
        25573 => X"B0",  -- 176
        25574 => X"AA",  -- 170
        25575 => X"AA",  -- 170
        25576 => X"B8",  -- 184
        25577 => X"BC",  -- 188
        25578 => X"B7",  -- 183
        25579 => X"AA",  -- 170
        25580 => X"A0",  -- 160
        25581 => X"A1",  -- 161
        25582 => X"A7",  -- 167
        25583 => X"A9",  -- 169
        25584 => X"A7",  -- 167
        25585 => X"B1",  -- 177
        25586 => X"BE",  -- 190
        25587 => X"C5",  -- 197
        25588 => X"CA",  -- 202
        25589 => X"CA",  -- 202
        25590 => X"C3",  -- 195
        25591 => X"BA",  -- 186
        25592 => X"B1",  -- 177
        25593 => X"A4",  -- 164
        25594 => X"9D",  -- 157
        25595 => X"A2",  -- 162
        25596 => X"A4",  -- 164
        25597 => X"A2",  -- 162
        25598 => X"A2",  -- 162
        25599 => X"A8",  -- 168
        25600 => X"6F",  -- 111
        25601 => X"6B",  -- 107
        25602 => X"67",  -- 103
        25603 => X"65",  -- 101
        25604 => X"67",  -- 103
        25605 => X"6C",  -- 108
        25606 => X"70",  -- 112
        25607 => X"73",  -- 115
        25608 => X"6F",  -- 111
        25609 => X"67",  -- 103
        25610 => X"5E",  -- 94
        25611 => X"5A",  -- 90
        25612 => X"5C",  -- 92
        25613 => X"61",  -- 97
        25614 => X"65",  -- 101
        25615 => X"66",  -- 102
        25616 => X"61",  -- 97
        25617 => X"61",  -- 97
        25618 => X"61",  -- 97
        25619 => X"61",  -- 97
        25620 => X"65",  -- 101
        25621 => X"6A",  -- 106
        25622 => X"69",  -- 105
        25623 => X"65",  -- 101
        25624 => X"64",  -- 100
        25625 => X"5A",  -- 90
        25626 => X"53",  -- 83
        25627 => X"57",  -- 87
        25628 => X"5D",  -- 93
        25629 => X"5E",  -- 94
        25630 => X"5C",  -- 92
        25631 => X"5A",  -- 90
        25632 => X"53",  -- 83
        25633 => X"32",  -- 50
        25634 => X"1D",  -- 29
        25635 => X"25",  -- 37
        25636 => X"30",  -- 48
        25637 => X"39",  -- 57
        25638 => X"4B",  -- 75
        25639 => X"63",  -- 99
        25640 => X"72",  -- 114
        25641 => X"8B",  -- 139
        25642 => X"A2",  -- 162
        25643 => X"A0",  -- 160
        25644 => X"89",  -- 137
        25645 => X"67",  -- 103
        25646 => X"46",  -- 70
        25647 => X"2F",  -- 47
        25648 => X"1D",  -- 29
        25649 => X"26",  -- 38
        25650 => X"40",  -- 64
        25651 => X"5B",  -- 91
        25652 => X"74",  -- 116
        25653 => X"69",  -- 105
        25654 => X"32",  -- 50
        25655 => X"12",  -- 18
        25656 => X"06",  -- 6
        25657 => X"04",  -- 4
        25658 => X"25",  -- 37
        25659 => X"5D",  -- 93
        25660 => X"7B",  -- 123
        25661 => X"91",  -- 145
        25662 => X"A7",  -- 167
        25663 => X"AE",  -- 174
        25664 => X"B6",  -- 182
        25665 => X"C4",  -- 196
        25666 => X"CD",  -- 205
        25667 => X"D4",  -- 212
        25668 => X"D0",  -- 208
        25669 => X"B2",  -- 178
        25670 => X"40",  -- 64
        25671 => X"07",  -- 7
        25672 => X"1D",  -- 29
        25673 => X"1C",  -- 28
        25674 => X"55",  -- 85
        25675 => X"6B",  -- 107
        25676 => X"7F",  -- 127
        25677 => X"AC",  -- 172
        25678 => X"9E",  -- 158
        25679 => X"8C",  -- 140
        25680 => X"8C",  -- 140
        25681 => X"7A",  -- 122
        25682 => X"7E",  -- 126
        25683 => X"77",  -- 119
        25684 => X"7C",  -- 124
        25685 => X"75",  -- 117
        25686 => X"89",  -- 137
        25687 => X"90",  -- 144
        25688 => X"8B",  -- 139
        25689 => X"87",  -- 135
        25690 => X"90",  -- 144
        25691 => X"75",  -- 117
        25692 => X"73",  -- 115
        25693 => X"5D",  -- 93
        25694 => X"1E",  -- 30
        25695 => X"2A",  -- 42
        25696 => X"65",  -- 101
        25697 => X"6E",  -- 110
        25698 => X"3F",  -- 63
        25699 => X"28",  -- 40
        25700 => X"20",  -- 32
        25701 => X"27",  -- 39
        25702 => X"3D",  -- 61
        25703 => X"6F",  -- 111
        25704 => X"7A",  -- 122
        25705 => X"7B",  -- 123
        25706 => X"8A",  -- 138
        25707 => X"89",  -- 137
        25708 => X"80",  -- 128
        25709 => X"85",  -- 133
        25710 => X"8D",  -- 141
        25711 => X"97",  -- 151
        25712 => X"9E",  -- 158
        25713 => X"AE",  -- 174
        25714 => X"C7",  -- 199
        25715 => X"C2",  -- 194
        25716 => X"8E",  -- 142
        25717 => X"95",  -- 149
        25718 => X"71",  -- 113
        25719 => X"20",  -- 32
        25720 => X"49",  -- 73
        25721 => X"8E",  -- 142
        25722 => X"CE",  -- 206
        25723 => X"DC",  -- 220
        25724 => X"D7",  -- 215
        25725 => X"DA",  -- 218
        25726 => X"D6",  -- 214
        25727 => X"CB",  -- 203
        25728 => X"C2",  -- 194
        25729 => X"BD",  -- 189
        25730 => X"AB",  -- 171
        25731 => X"9E",  -- 158
        25732 => X"83",  -- 131
        25733 => X"3C",  -- 60
        25734 => X"0B",  -- 11
        25735 => X"12",  -- 18
        25736 => X"0F",  -- 15
        25737 => X"32",  -- 50
        25738 => X"6F",  -- 111
        25739 => X"92",  -- 146
        25740 => X"8B",  -- 139
        25741 => X"83",  -- 131
        25742 => X"77",  -- 119
        25743 => X"5F",  -- 95
        25744 => X"4A",  -- 74
        25745 => X"35",  -- 53
        25746 => X"25",  -- 37
        25747 => X"34",  -- 52
        25748 => X"55",  -- 85
        25749 => X"70",  -- 112
        25750 => X"8F",  -- 143
        25751 => X"B0",  -- 176
        25752 => X"BA",  -- 186
        25753 => X"AA",  -- 170
        25754 => X"A5",  -- 165
        25755 => X"AE",  -- 174
        25756 => X"8E",  -- 142
        25757 => X"60",  -- 96
        25758 => X"50",  -- 80
        25759 => X"3E",  -- 62
        25760 => X"56",  -- 86
        25761 => X"52",  -- 82
        25762 => X"29",  -- 41
        25763 => X"34",  -- 52
        25764 => X"82",  -- 130
        25765 => X"A8",  -- 168
        25766 => X"97",  -- 151
        25767 => X"74",  -- 116
        25768 => X"71",  -- 113
        25769 => X"5E",  -- 94
        25770 => X"75",  -- 117
        25771 => X"98",  -- 152
        25772 => X"9A",  -- 154
        25773 => X"90",  -- 144
        25774 => X"7F",  -- 127
        25775 => X"60",  -- 96
        25776 => X"70",  -- 112
        25777 => X"7F",  -- 127
        25778 => X"91",  -- 145
        25779 => X"9B",  -- 155
        25780 => X"94",  -- 148
        25781 => X"84",  -- 132
        25782 => X"71",  -- 113
        25783 => X"65",  -- 101
        25784 => X"53",  -- 83
        25785 => X"43",  -- 67
        25786 => X"31",  -- 49
        25787 => X"22",  -- 34
        25788 => X"16",  -- 22
        25789 => X"13",  -- 19
        25790 => X"1F",  -- 31
        25791 => X"2F",  -- 47
        25792 => X"5A",  -- 90
        25793 => X"6C",  -- 108
        25794 => X"93",  -- 147
        25795 => X"98",  -- 152
        25796 => X"96",  -- 150
        25797 => X"AB",  -- 171
        25798 => X"AF",  -- 175
        25799 => X"A8",  -- 168
        25800 => X"A8",  -- 168
        25801 => X"AE",  -- 174
        25802 => X"B5",  -- 181
        25803 => X"BB",  -- 187
        25804 => X"B8",  -- 184
        25805 => X"B2",  -- 178
        25806 => X"AB",  -- 171
        25807 => X"A8",  -- 168
        25808 => X"C1",  -- 193
        25809 => X"C6",  -- 198
        25810 => X"C5",  -- 197
        25811 => X"BE",  -- 190
        25812 => X"BC",  -- 188
        25813 => X"BC",  -- 188
        25814 => X"BB",  -- 187
        25815 => X"B9",  -- 185
        25816 => X"B9",  -- 185
        25817 => X"BD",  -- 189
        25818 => X"C2",  -- 194
        25819 => X"C7",  -- 199
        25820 => X"C9",  -- 201
        25821 => X"C8",  -- 200
        25822 => X"C7",  -- 199
        25823 => X"C6",  -- 198
        25824 => X"B0",  -- 176
        25825 => X"A3",  -- 163
        25826 => X"94",  -- 148
        25827 => X"92",  -- 146
        25828 => X"99",  -- 153
        25829 => X"A5",  -- 165
        25830 => X"B1",  -- 177
        25831 => X"B9",  -- 185
        25832 => X"AE",  -- 174
        25833 => X"B0",  -- 176
        25834 => X"B0",  -- 176
        25835 => X"B0",  -- 176
        25836 => X"B1",  -- 177
        25837 => X"B2",  -- 178
        25838 => X"AC",  -- 172
        25839 => X"A5",  -- 165
        25840 => X"9E",  -- 158
        25841 => X"95",  -- 149
        25842 => X"8F",  -- 143
        25843 => X"95",  -- 149
        25844 => X"94",  -- 148
        25845 => X"80",  -- 128
        25846 => X"60",  -- 96
        25847 => X"46",  -- 70
        25848 => X"37",  -- 55
        25849 => X"35",  -- 53
        25850 => X"39",  -- 57
        25851 => X"4E",  -- 78
        25852 => X"73",  -- 115
        25853 => X"92",  -- 146
        25854 => X"96",  -- 150
        25855 => X"8C",  -- 140
        25856 => X"93",  -- 147
        25857 => X"9E",  -- 158
        25858 => X"A4",  -- 164
        25859 => X"AA",  -- 170
        25860 => X"B4",  -- 180
        25861 => X"B9",  -- 185
        25862 => X"C2",  -- 194
        25863 => X"CF",  -- 207
        25864 => X"D0",  -- 208
        25865 => X"CC",  -- 204
        25866 => X"CE",  -- 206
        25867 => X"CB",  -- 203
        25868 => X"C2",  -- 194
        25869 => X"C5",  -- 197
        25870 => X"B1",  -- 177
        25871 => X"88",  -- 136
        25872 => X"4C",  -- 76
        25873 => X"19",  -- 25
        25874 => X"26",  -- 38
        25875 => X"64",  -- 100
        25876 => X"77",  -- 119
        25877 => X"79",  -- 121
        25878 => X"8F",  -- 143
        25879 => X"A5",  -- 165
        25880 => X"9A",  -- 154
        25881 => X"92",  -- 146
        25882 => X"7F",  -- 127
        25883 => X"98",  -- 152
        25884 => X"A2",  -- 162
        25885 => X"A0",  -- 160
        25886 => X"8B",  -- 139
        25887 => X"9D",  -- 157
        25888 => X"98",  -- 152
        25889 => X"9D",  -- 157
        25890 => X"AB",  -- 171
        25891 => X"B3",  -- 179
        25892 => X"AD",  -- 173
        25893 => X"AB",  -- 171
        25894 => X"AC",  -- 172
        25895 => X"A6",  -- 166
        25896 => X"B0",  -- 176
        25897 => X"B3",  -- 179
        25898 => X"AE",  -- 174
        25899 => X"A3",  -- 163
        25900 => X"9F",  -- 159
        25901 => X"A5",  -- 165
        25902 => X"AA",  -- 170
        25903 => X"AB",  -- 171
        25904 => X"A6",  -- 166
        25905 => X"B2",  -- 178
        25906 => X"BA",  -- 186
        25907 => X"BF",  -- 191
        25908 => X"C6",  -- 198
        25909 => X"CB",  -- 203
        25910 => X"C4",  -- 196
        25911 => X"B7",  -- 183
        25912 => X"AE",  -- 174
        25913 => X"A5",  -- 165
        25914 => X"A1",  -- 161
        25915 => X"A5",  -- 165
        25916 => X"A9",  -- 169
        25917 => X"A5",  -- 165
        25918 => X"A1",  -- 161
        25919 => X"A1",  -- 161
        25920 => X"69",  -- 105
        25921 => X"67",  -- 103
        25922 => X"65",  -- 101
        25923 => X"64",  -- 100
        25924 => X"65",  -- 101
        25925 => X"66",  -- 102
        25926 => X"66",  -- 102
        25927 => X"66",  -- 102
        25928 => X"6E",  -- 110
        25929 => X"68",  -- 104
        25930 => X"61",  -- 97
        25931 => X"5D",  -- 93
        25932 => X"5D",  -- 93
        25933 => X"60",  -- 96
        25934 => X"64",  -- 100
        25935 => X"67",  -- 103
        25936 => X"68",  -- 104
        25937 => X"6C",  -- 108
        25938 => X"6D",  -- 109
        25939 => X"6E",  -- 110
        25940 => X"71",  -- 113
        25941 => X"74",  -- 116
        25942 => X"72",  -- 114
        25943 => X"6E",  -- 110
        25944 => X"65",  -- 101
        25945 => X"5D",  -- 93
        25946 => X"56",  -- 86
        25947 => X"58",  -- 88
        25948 => X"5D",  -- 93
        25949 => X"5D",  -- 93
        25950 => X"5C",  -- 92
        25951 => X"5D",  -- 93
        25952 => X"4E",  -- 78
        25953 => X"2A",  -- 42
        25954 => X"13",  -- 19
        25955 => X"19",  -- 25
        25956 => X"26",  -- 38
        25957 => X"2F",  -- 47
        25958 => X"47",  -- 71
        25959 => X"64",  -- 100
        25960 => X"86",  -- 134
        25961 => X"95",  -- 149
        25962 => X"9C",  -- 156
        25963 => X"8D",  -- 141
        25964 => X"6E",  -- 110
        25965 => X"4D",  -- 77
        25966 => X"31",  -- 49
        25967 => X"1F",  -- 31
        25968 => X"18",  -- 24
        25969 => X"35",  -- 53
        25970 => X"5C",  -- 92
        25971 => X"6B",  -- 107
        25972 => X"6C",  -- 108
        25973 => X"55",  -- 85
        25974 => X"26",  -- 38
        25975 => X"13",  -- 19
        25976 => X"09",  -- 9
        25977 => X"0A",  -- 10
        25978 => X"31",  -- 49
        25979 => X"6B",  -- 107
        25980 => X"90",  -- 144
        25981 => X"A2",  -- 162
        25982 => X"AD",  -- 173
        25983 => X"AC",  -- 172
        25984 => X"BC",  -- 188
        25985 => X"C7",  -- 199
        25986 => X"CD",  -- 205
        25987 => X"CF",  -- 207
        25988 => X"C6",  -- 198
        25989 => X"B8",  -- 184
        25990 => X"77",  -- 119
        25991 => X"63",  -- 99
        25992 => X"60",  -- 96
        25993 => X"7D",  -- 125
        25994 => X"B4",  -- 180
        25995 => X"CA",  -- 202
        25996 => X"C3",  -- 195
        25997 => X"BB",  -- 187
        25998 => X"A6",  -- 166
        25999 => X"8D",  -- 141
        26000 => X"7D",  -- 125
        26001 => X"7D",  -- 125
        26002 => X"6A",  -- 106
        26003 => X"61",  -- 97
        26004 => X"6F",  -- 111
        26005 => X"86",  -- 134
        26006 => X"8C",  -- 140
        26007 => X"8D",  -- 141
        26008 => X"93",  -- 147
        26009 => X"84",  -- 132
        26010 => X"7C",  -- 124
        26011 => X"6D",  -- 109
        26012 => X"45",  -- 69
        26013 => X"4A",  -- 74
        26014 => X"28",  -- 40
        26015 => X"34",  -- 52
        26016 => X"6F",  -- 111
        26017 => X"6C",  -- 108
        26018 => X"3C",  -- 60
        26019 => X"25",  -- 37
        26020 => X"20",  -- 32
        26021 => X"31",  -- 49
        26022 => X"44",  -- 68
        26023 => X"67",  -- 103
        26024 => X"6C",  -- 108
        26025 => X"62",  -- 98
        26026 => X"6C",  -- 108
        26027 => X"70",  -- 112
        26028 => X"65",  -- 101
        26029 => X"56",  -- 86
        26030 => X"56",  -- 86
        26031 => X"61",  -- 97
        26032 => X"72",  -- 114
        26033 => X"8D",  -- 141
        26034 => X"B7",  -- 183
        26035 => X"DD",  -- 221
        26036 => X"D1",  -- 209
        26037 => X"D0",  -- 208
        26038 => X"B7",  -- 183
        26039 => X"97",  -- 151
        26040 => X"A3",  -- 163
        26041 => X"C4",  -- 196
        26042 => X"DD",  -- 221
        26043 => X"DF",  -- 223
        26044 => X"DE",  -- 222
        26045 => X"E1",  -- 225
        26046 => X"DA",  -- 218
        26047 => X"C9",  -- 201
        26048 => X"CE",  -- 206
        26049 => X"BE",  -- 190
        26050 => X"B8",  -- 184
        26051 => X"A1",  -- 161
        26052 => X"75",  -- 117
        26053 => X"59",  -- 89
        26054 => X"39",  -- 57
        26055 => X"0A",  -- 10
        26056 => X"0C",  -- 12
        26057 => X"2B",  -- 43
        26058 => X"6B",  -- 107
        26059 => X"9D",  -- 157
        26060 => X"A2",  -- 162
        26061 => X"94",  -- 148
        26062 => X"82",  -- 130
        26063 => X"70",  -- 112
        26064 => X"56",  -- 86
        26065 => X"4C",  -- 76
        26066 => X"37",  -- 55
        26067 => X"31",  -- 49
        26068 => X"3F",  -- 63
        26069 => X"57",  -- 87
        26070 => X"79",  -- 121
        26071 => X"9B",  -- 155
        26072 => X"B8",  -- 184
        26073 => X"B9",  -- 185
        26074 => X"AA",  -- 170
        26075 => X"94",  -- 148
        26076 => X"74",  -- 116
        26077 => X"62",  -- 98
        26078 => X"56",  -- 86
        26079 => X"32",  -- 50
        26080 => X"27",  -- 39
        26081 => X"28",  -- 40
        26082 => X"36",  -- 54
        26083 => X"6A",  -- 106
        26084 => X"99",  -- 153
        26085 => X"AF",  -- 175
        26086 => X"AA",  -- 170
        26087 => X"88",  -- 136
        26088 => X"77",  -- 119
        26089 => X"63",  -- 99
        26090 => X"6C",  -- 108
        26091 => X"85",  -- 133
        26092 => X"8D",  -- 141
        26093 => X"95",  -- 149
        26094 => X"8E",  -- 142
        26095 => X"6F",  -- 111
        26096 => X"68",  -- 104
        26097 => X"72",  -- 114
        26098 => X"81",  -- 129
        26099 => X"8A",  -- 138
        26100 => X"88",  -- 136
        26101 => X"7E",  -- 126
        26102 => X"72",  -- 114
        26103 => X"69",  -- 105
        26104 => X"5E",  -- 94
        26105 => X"52",  -- 82
        26106 => X"40",  -- 64
        26107 => X"2C",  -- 44
        26108 => X"19",  -- 25
        26109 => X"12",  -- 18
        26110 => X"20",  -- 32
        26111 => X"33",  -- 51
        26112 => X"55",  -- 85
        26113 => X"5C",  -- 92
        26114 => X"7C",  -- 124
        26115 => X"8C",  -- 140
        26116 => X"9B",  -- 155
        26117 => X"B1",  -- 177
        26118 => X"B0",  -- 176
        26119 => X"AE",  -- 174
        26120 => X"AA",  -- 170
        26121 => X"AC",  -- 172
        26122 => X"B4",  -- 180
        26123 => X"BF",  -- 191
        26124 => X"C6",  -- 198
        26125 => X"C5",  -- 197
        26126 => X"BB",  -- 187
        26127 => X"B2",  -- 178
        26128 => X"B1",  -- 177
        26129 => X"B6",  -- 182
        26130 => X"BA",  -- 186
        26131 => X"BA",  -- 186
        26132 => X"BD",  -- 189
        26133 => X"C1",  -- 193
        26134 => X"C2",  -- 194
        26135 => X"BF",  -- 191
        26136 => X"BB",  -- 187
        26137 => X"BC",  -- 188
        26138 => X"C1",  -- 193
        26139 => X"C4",  -- 196
        26140 => X"C6",  -- 198
        26141 => X"C5",  -- 197
        26142 => X"C2",  -- 194
        26143 => X"C0",  -- 192
        26144 => X"A7",  -- 167
        26145 => X"8C",  -- 140
        26146 => X"75",  -- 117
        26147 => X"79",  -- 121
        26148 => X"93",  -- 147
        26149 => X"AD",  -- 173
        26150 => X"BA",  -- 186
        26151 => X"BD",  -- 189
        26152 => X"B8",  -- 184
        26153 => X"BC",  -- 188
        26154 => X"BD",  -- 189
        26155 => X"B9",  -- 185
        26156 => X"B5",  -- 181
        26157 => X"B2",  -- 178
        26158 => X"AD",  -- 173
        26159 => X"A8",  -- 168
        26160 => X"9D",  -- 157
        26161 => X"9B",  -- 155
        26162 => X"97",  -- 151
        26163 => X"8D",  -- 141
        26164 => X"79",  -- 121
        26165 => X"64",  -- 100
        26166 => X"55",  -- 85
        26167 => X"52",  -- 82
        26168 => X"45",  -- 69
        26169 => X"2A",  -- 42
        26170 => X"28",  -- 40
        26171 => X"4B",  -- 75
        26172 => X"72",  -- 114
        26173 => X"86",  -- 134
        26174 => X"99",  -- 153
        26175 => X"AE",  -- 174
        26176 => X"A9",  -- 169
        26177 => X"B1",  -- 177
        26178 => X"B2",  -- 178
        26179 => X"B2",  -- 178
        26180 => X"BA",  -- 186
        26181 => X"BD",  -- 189
        26182 => X"C0",  -- 192
        26183 => X"CA",  -- 202
        26184 => X"CE",  -- 206
        26185 => X"CB",  -- 203
        26186 => X"CE",  -- 206
        26187 => X"CB",  -- 203
        26188 => X"C8",  -- 200
        26189 => X"C6",  -- 198
        26190 => X"A9",  -- 169
        26191 => X"78",  -- 120
        26192 => X"31",  -- 49
        26193 => X"1A",  -- 26
        26194 => X"2C",  -- 44
        26195 => X"5D",  -- 93
        26196 => X"7F",  -- 127
        26197 => X"99",  -- 153
        26198 => X"A4",  -- 164
        26199 => X"99",  -- 153
        26200 => X"A7",  -- 167
        26201 => X"AC",  -- 172
        26202 => X"A0",  -- 160
        26203 => X"92",  -- 146
        26204 => X"A0",  -- 160
        26205 => X"9E",  -- 158
        26206 => X"96",  -- 150
        26207 => X"98",  -- 152
        26208 => X"9A",  -- 154
        26209 => X"9D",  -- 157
        26210 => X"AA",  -- 170
        26211 => X"B0",  -- 176
        26212 => X"AC",  -- 172
        26213 => X"AA",  -- 170
        26214 => X"AB",  -- 171
        26215 => X"A7",  -- 167
        26216 => X"AC",  -- 172
        26217 => X"A9",  -- 169
        26218 => X"A2",  -- 162
        26219 => X"99",  -- 153
        26220 => X"9A",  -- 154
        26221 => X"A3",  -- 163
        26222 => X"A7",  -- 167
        26223 => X"A6",  -- 166
        26224 => X"AE",  -- 174
        26225 => X"B2",  -- 178
        26226 => X"B9",  -- 185
        26227 => X"C0",  -- 192
        26228 => X"C8",  -- 200
        26229 => X"CD",  -- 205
        26230 => X"C6",  -- 198
        26231 => X"BD",  -- 189
        26232 => X"B4",  -- 180
        26233 => X"AA",  -- 170
        26234 => X"A1",  -- 161
        26235 => X"A0",  -- 160
        26236 => X"A0",  -- 160
        26237 => X"9F",  -- 159
        26238 => X"9F",  -- 159
        26239 => X"A2",  -- 162
        26240 => X"6B",  -- 107
        26241 => X"6B",  -- 107
        26242 => X"6A",  -- 106
        26243 => X"6A",  -- 106
        26244 => X"69",  -- 105
        26245 => X"66",  -- 102
        26246 => X"63",  -- 99
        26247 => X"60",  -- 96
        26248 => X"67",  -- 103
        26249 => X"64",  -- 100
        26250 => X"60",  -- 96
        26251 => X"5D",  -- 93
        26252 => X"5C",  -- 92
        26253 => X"60",  -- 96
        26254 => X"66",  -- 102
        26255 => X"6B",  -- 107
        26256 => X"74",  -- 116
        26257 => X"7C",  -- 124
        26258 => X"83",  -- 131
        26259 => X"85",  -- 133
        26260 => X"86",  -- 134
        26261 => X"86",  -- 134
        26262 => X"84",  -- 132
        26263 => X"80",  -- 128
        26264 => X"72",  -- 114
        26265 => X"69",  -- 105
        26266 => X"61",  -- 97
        26267 => X"60",  -- 96
        26268 => X"60",  -- 96
        26269 => X"5E",  -- 94
        26270 => X"5B",  -- 91
        26271 => X"5A",  -- 90
        26272 => X"5A",  -- 90
        26273 => X"41",  -- 65
        26274 => X"2D",  -- 45
        26275 => X"28",  -- 40
        26276 => X"29",  -- 41
        26277 => X"34",  -- 52
        26278 => X"58",  -- 88
        26279 => X"7F",  -- 127
        26280 => X"A0",  -- 160
        26281 => X"A0",  -- 160
        26282 => X"95",  -- 149
        26283 => X"79",  -- 121
        26284 => X"55",  -- 85
        26285 => X"39",  -- 57
        26286 => X"2A",  -- 42
        26287 => X"25",  -- 37
        26288 => X"24",  -- 36
        26289 => X"42",  -- 66
        26290 => X"6A",  -- 106
        26291 => X"75",  -- 117
        26292 => X"6F",  -- 111
        26293 => X"4E",  -- 78
        26294 => X"1C",  -- 28
        26295 => X"09",  -- 9
        26296 => X"0E",  -- 14
        26297 => X"1C",  -- 28
        26298 => X"46",  -- 70
        26299 => X"78",  -- 120
        26300 => X"95",  -- 149
        26301 => X"A8",  -- 168
        26302 => X"B7",  -- 183
        26303 => X"BC",  -- 188
        26304 => X"C4",  -- 196
        26305 => X"C8",  -- 200
        26306 => X"CB",  -- 203
        26307 => X"CF",  -- 207
        26308 => X"CC",  -- 204
        26309 => X"C9",  -- 201
        26310 => X"B5",  -- 181
        26311 => X"C1",  -- 193
        26312 => X"CA",  -- 202
        26313 => X"C9",  -- 201
        26314 => X"C9",  -- 201
        26315 => X"D9",  -- 217
        26316 => X"C3",  -- 195
        26317 => X"8E",  -- 142
        26318 => X"73",  -- 115
        26319 => X"66",  -- 102
        26320 => X"3C",  -- 60
        26321 => X"35",  -- 53
        26322 => X"3D",  -- 61
        26323 => X"71",  -- 113
        26324 => X"80",  -- 128
        26325 => X"94",  -- 148
        26326 => X"88",  -- 136
        26327 => X"82",  -- 130
        26328 => X"75",  -- 117
        26329 => X"64",  -- 100
        26330 => X"35",  -- 53
        26331 => X"2E",  -- 46
        26332 => X"39",  -- 57
        26333 => X"31",  -- 49
        26334 => X"22",  -- 34
        26335 => X"45",  -- 69
        26336 => X"68",  -- 104
        26337 => X"70",  -- 112
        26338 => X"5B",  -- 91
        26339 => X"3E",  -- 62
        26340 => X"1B",  -- 27
        26341 => X"20",  -- 32
        26342 => X"34",  -- 52
        26343 => X"56",  -- 86
        26344 => X"75",  -- 117
        26345 => X"5A",  -- 90
        26346 => X"36",  -- 54
        26347 => X"20",  -- 32
        26348 => X"14",  -- 20
        26349 => X"0F",  -- 15
        26350 => X"11",  -- 17
        26351 => X"17",  -- 23
        26352 => X"26",  -- 38
        26353 => X"2B",  -- 43
        26354 => X"54",  -- 84
        26355 => X"B6",  -- 182
        26356 => X"E4",  -- 228
        26357 => X"E2",  -- 226
        26358 => X"CD",  -- 205
        26359 => X"DE",  -- 222
        26360 => X"E0",  -- 224
        26361 => X"E4",  -- 228
        26362 => X"E2",  -- 226
        26363 => X"DE",  -- 222
        26364 => X"E1",  -- 225
        26365 => X"E6",  -- 230
        26366 => X"DE",  -- 222
        26367 => X"D0",  -- 208
        26368 => X"CB",  -- 203
        26369 => X"D2",  -- 210
        26370 => X"BB",  -- 187
        26371 => X"9B",  -- 155
        26372 => X"95",  -- 149
        26373 => X"89",  -- 137
        26374 => X"55",  -- 85
        26375 => X"20",  -- 32
        26376 => X"3A",  -- 58
        26377 => X"40",  -- 64
        26378 => X"62",  -- 98
        26379 => X"8F",  -- 143
        26380 => X"9E",  -- 158
        26381 => X"9A",  -- 154
        26382 => X"96",  -- 150
        26383 => X"92",  -- 146
        26384 => X"64",  -- 100
        26385 => X"60",  -- 96
        26386 => X"49",  -- 73
        26387 => X"2E",  -- 46
        26388 => X"28",  -- 40
        26389 => X"38",  -- 56
        26390 => X"59",  -- 89
        26391 => X"7B",  -- 123
        26392 => X"9C",  -- 156
        26393 => X"B5",  -- 181
        26394 => X"BF",  -- 191
        26395 => X"AA",  -- 170
        26396 => X"75",  -- 117
        26397 => X"4C",  -- 76
        26398 => X"45",  -- 69
        26399 => X"38",  -- 56
        26400 => X"1C",  -- 28
        26401 => X"14",  -- 20
        26402 => X"47",  -- 71
        26403 => X"9A",  -- 154
        26404 => X"B1",  -- 177
        26405 => X"B1",  -- 177
        26406 => X"B4",  -- 180
        26407 => X"91",  -- 145
        26408 => X"82",  -- 130
        26409 => X"6E",  -- 110
        26410 => X"6A",  -- 106
        26411 => X"75",  -- 117
        26412 => X"7F",  -- 127
        26413 => X"91",  -- 145
        26414 => X"8D",  -- 141
        26415 => X"6F",  -- 111
        26416 => X"71",  -- 113
        26417 => X"76",  -- 118
        26418 => X"7D",  -- 125
        26419 => X"81",  -- 129
        26420 => X"7F",  -- 127
        26421 => X"78",  -- 120
        26422 => X"6F",  -- 111
        26423 => X"69",  -- 105
        26424 => X"63",  -- 99
        26425 => X"58",  -- 88
        26426 => X"49",  -- 73
        26427 => X"31",  -- 49
        26428 => X"18",  -- 24
        26429 => X"0F",  -- 15
        26430 => X"1F",  -- 31
        26431 => X"38",  -- 56
        26432 => X"63",  -- 99
        26433 => X"64",  -- 100
        26434 => X"70",  -- 112
        26435 => X"7A",  -- 122
        26436 => X"92",  -- 146
        26437 => X"A3",  -- 163
        26438 => X"A2",  -- 162
        26439 => X"AE",  -- 174
        26440 => X"AF",  -- 175
        26441 => X"AE",  -- 174
        26442 => X"B1",  -- 177
        26443 => X"BD",  -- 189
        26444 => X"CB",  -- 203
        26445 => X"D0",  -- 208
        26446 => X"CA",  -- 202
        26447 => X"C1",  -- 193
        26448 => X"C3",  -- 195
        26449 => X"C5",  -- 197
        26450 => X"C5",  -- 197
        26451 => X"C4",  -- 196
        26452 => X"C3",  -- 195
        26453 => X"C2",  -- 194
        26454 => X"BF",  -- 191
        26455 => X"B9",  -- 185
        26456 => X"BB",  -- 187
        26457 => X"BC",  -- 188
        26458 => X"BF",  -- 191
        26459 => X"C3",  -- 195
        26460 => X"C8",  -- 200
        26461 => X"CB",  -- 203
        26462 => X"C9",  -- 201
        26463 => X"C7",  -- 199
        26464 => X"AE",  -- 174
        26465 => X"8E",  -- 142
        26466 => X"74",  -- 116
        26467 => X"78",  -- 120
        26468 => X"92",  -- 146
        26469 => X"A8",  -- 168
        26470 => X"B1",  -- 177
        26471 => X"B2",  -- 178
        26472 => X"B7",  -- 183
        26473 => X"BD",  -- 189
        26474 => X"BE",  -- 190
        26475 => X"BA",  -- 186
        26476 => X"B2",  -- 178
        26477 => X"AF",  -- 175
        26478 => X"AD",  -- 173
        26479 => X"AB",  -- 171
        26480 => X"99",  -- 153
        26481 => X"94",  -- 148
        26482 => X"8E",  -- 142
        26483 => X"8C",  -- 140
        26484 => X"83",  -- 131
        26485 => X"70",  -- 112
        26486 => X"5A",  -- 90
        26487 => X"4C",  -- 76
        26488 => X"4B",  -- 75
        26489 => X"31",  -- 49
        26490 => X"31",  -- 49
        26491 => X"57",  -- 87
        26492 => X"75",  -- 117
        26493 => X"7B",  -- 123
        26494 => X"8A",  -- 138
        26495 => X"A2",  -- 162
        26496 => X"AE",  -- 174
        26497 => X"B5",  -- 181
        26498 => X"B5",  -- 181
        26499 => X"B7",  -- 183
        26500 => X"C2",  -- 194
        26501 => X"C5",  -- 197
        26502 => X"C6",  -- 198
        26503 => X"CD",  -- 205
        26504 => X"C3",  -- 195
        26505 => X"C4",  -- 196
        26506 => X"C7",  -- 199
        26507 => X"C9",  -- 201
        26508 => X"CB",  -- 203
        26509 => X"C5",  -- 197
        26510 => X"9B",  -- 155
        26511 => X"63",  -- 99
        26512 => X"26",  -- 38
        26513 => X"27",  -- 39
        26514 => X"47",  -- 71
        26515 => X"71",  -- 113
        26516 => X"91",  -- 145
        26517 => X"AB",  -- 171
        26518 => X"AF",  -- 175
        26519 => X"9C",  -- 156
        26520 => X"90",  -- 144
        26521 => X"A8",  -- 168
        26522 => X"AA",  -- 170
        26523 => X"89",  -- 137
        26524 => X"9F",  -- 159
        26525 => X"A2",  -- 162
        26526 => X"A8",  -- 168
        26527 => X"9C",  -- 156
        26528 => X"98",  -- 152
        26529 => X"99",  -- 153
        26530 => X"A2",  -- 162
        26531 => X"A7",  -- 167
        26532 => X"A3",  -- 163
        26533 => X"A3",  -- 163
        26534 => X"A7",  -- 167
        26535 => X"A2",  -- 162
        26536 => X"A9",  -- 169
        26537 => X"A0",  -- 160
        26538 => X"95",  -- 149
        26539 => X"92",  -- 146
        26540 => X"99",  -- 153
        26541 => X"A3",  -- 163
        26542 => X"A7",  -- 167
        26543 => X"A7",  -- 167
        26544 => X"B1",  -- 177
        26545 => X"AD",  -- 173
        26546 => X"B0",  -- 176
        26547 => X"BE",  -- 190
        26548 => X"C9",  -- 201
        26549 => X"CB",  -- 203
        26550 => X"C4",  -- 196
        26551 => X"BF",  -- 191
        26552 => X"C3",  -- 195
        26553 => X"BB",  -- 187
        26554 => X"AF",  -- 175
        26555 => X"A7",  -- 167
        26556 => X"A1",  -- 161
        26557 => X"9A",  -- 154
        26558 => X"97",  -- 151
        26559 => X"96",  -- 150
        26560 => X"6E",  -- 110
        26561 => X"6E",  -- 110
        26562 => X"6F",  -- 111
        26563 => X"6F",  -- 111
        26564 => X"6E",  -- 110
        26565 => X"6A",  -- 106
        26566 => X"66",  -- 102
        26567 => X"62",  -- 98
        26568 => X"60",  -- 96
        26569 => X"60",  -- 96
        26570 => X"60",  -- 96
        26571 => X"5E",  -- 94
        26572 => X"5F",  -- 95
        26573 => X"63",  -- 99
        26574 => X"6B",  -- 107
        26575 => X"73",  -- 115
        26576 => X"7F",  -- 127
        26577 => X"89",  -- 137
        26578 => X"94",  -- 148
        26579 => X"98",  -- 152
        26580 => X"98",  -- 152
        26581 => X"97",  -- 151
        26582 => X"94",  -- 148
        26583 => X"91",  -- 145
        26584 => X"82",  -- 130
        26585 => X"7A",  -- 122
        26586 => X"72",  -- 114
        26587 => X"6D",  -- 109
        26588 => X"67",  -- 103
        26589 => X"5E",  -- 94
        26590 => X"56",  -- 86
        26591 => X"55",  -- 85
        26592 => X"52",  -- 82
        26593 => X"50",  -- 80
        26594 => X"45",  -- 69
        26595 => X"31",  -- 49
        26596 => X"28",  -- 40
        26597 => X"3E",  -- 62
        26598 => X"6F",  -- 111
        26599 => X"97",  -- 151
        26600 => X"A2",  -- 162
        26601 => X"94",  -- 148
        26602 => X"7D",  -- 125
        26603 => X"5D",  -- 93
        26604 => X"3E",  -- 62
        26605 => X"31",  -- 49
        26606 => X"36",  -- 54
        26607 => X"3F",  -- 63
        26608 => X"5F",  -- 95
        26609 => X"62",  -- 98
        26610 => X"74",  -- 116
        26611 => X"80",  -- 128
        26612 => X"7D",  -- 125
        26613 => X"54",  -- 84
        26614 => X"18",  -- 24
        26615 => X"03",  -- 3
        26616 => X"04",  -- 4
        26617 => X"28",  -- 40
        26618 => X"60",  -- 96
        26619 => X"88",  -- 136
        26620 => X"9A",  -- 154
        26621 => X"AC",  -- 172
        26622 => X"C1",  -- 193
        26623 => X"D0",  -- 208
        26624 => X"CE",  -- 206
        26625 => X"CB",  -- 203
        26626 => X"CC",  -- 204
        26627 => X"D4",  -- 212
        26628 => X"D6",  -- 214
        26629 => X"D3",  -- 211
        26630 => X"CD",  -- 205
        26631 => X"D8",  -- 216
        26632 => X"CB",  -- 203
        26633 => X"D7",  -- 215
        26634 => X"D1",  -- 209
        26635 => X"B1",  -- 177
        26636 => X"73",  -- 115
        26637 => X"30",  -- 48
        26638 => X"11",  -- 17
        26639 => X"13",  -- 19
        26640 => X"0E",  -- 14
        26641 => X"0A",  -- 10
        26642 => X"34",  -- 52
        26643 => X"80",  -- 128
        26644 => X"84",  -- 132
        26645 => X"8D",  -- 141
        26646 => X"84",  -- 132
        26647 => X"63",  -- 99
        26648 => X"32",  -- 50
        26649 => X"22",  -- 34
        26650 => X"19",  -- 25
        26651 => X"1E",  -- 30
        26652 => X"47",  -- 71
        26653 => X"18",  -- 24
        26654 => X"32",  -- 50
        26655 => X"55",  -- 85
        26656 => X"5F",  -- 95
        26657 => X"6D",  -- 109
        26658 => X"80",  -- 128
        26659 => X"75",  -- 117
        26660 => X"3D",  -- 61
        26661 => X"2D",  -- 45
        26662 => X"2D",  -- 45
        26663 => X"45",  -- 69
        26664 => X"5D",  -- 93
        26665 => X"62",  -- 98
        26666 => X"41",  -- 65
        26667 => X"18",  -- 24
        26668 => X"06",  -- 6
        26669 => X"09",  -- 9
        26670 => X"0F",  -- 15
        26671 => X"07",  -- 7
        26672 => X"0A",  -- 10
        26673 => X"05",  -- 5
        26674 => X"16",  -- 22
        26675 => X"69",  -- 105
        26676 => X"B4",  -- 180
        26677 => X"E4",  -- 228
        26678 => X"E1",  -- 225
        26679 => X"E3",  -- 227
        26680 => X"E4",  -- 228
        26681 => X"E4",  -- 228
        26682 => X"E1",  -- 225
        26683 => X"E0",  -- 224
        26684 => X"E1",  -- 225
        26685 => X"E2",  -- 226
        26686 => X"E0",  -- 224
        26687 => X"DC",  -- 220
        26688 => X"CE",  -- 206
        26689 => X"D0",  -- 208
        26690 => X"B9",  -- 185
        26691 => X"AA",  -- 170
        26692 => X"B5",  -- 181
        26693 => X"9E",  -- 158
        26694 => X"5C",  -- 92
        26695 => X"2E",  -- 46
        26696 => X"16",  -- 22
        26697 => X"1E",  -- 30
        26698 => X"42",  -- 66
        26699 => X"79",  -- 121
        26700 => X"9E",  -- 158
        26701 => X"A5",  -- 165
        26702 => X"9D",  -- 157
        26703 => X"97",  -- 151
        26704 => X"7D",  -- 125
        26705 => X"76",  -- 118
        26706 => X"5D",  -- 93
        26707 => X"3F",  -- 63
        26708 => X"31",  -- 49
        26709 => X"33",  -- 51
        26710 => X"4A",  -- 74
        26711 => X"66",  -- 102
        26712 => X"98",  -- 152
        26713 => X"B0",  -- 176
        26714 => X"BE",  -- 190
        26715 => X"C6",  -- 198
        26716 => X"AE",  -- 174
        26717 => X"87",  -- 135
        26718 => X"6A",  -- 106
        26719 => X"4B",  -- 75
        26720 => X"40",  -- 64
        26721 => X"28",  -- 40
        26722 => X"4F",  -- 79
        26723 => X"9F",  -- 159
        26724 => X"B8",  -- 184
        26725 => X"B4",  -- 180
        26726 => X"B5",  -- 181
        26727 => X"93",  -- 147
        26728 => X"6C",  -- 108
        26729 => X"5C",  -- 92
        26730 => X"5A",  -- 90
        26731 => X"6C",  -- 108
        26732 => X"7E",  -- 126
        26733 => X"91",  -- 145
        26734 => X"90",  -- 144
        26735 => X"7D",  -- 125
        26736 => X"77",  -- 119
        26737 => X"7A",  -- 122
        26738 => X"7C",  -- 124
        26739 => X"7F",  -- 127
        26740 => X"7C",  -- 124
        26741 => X"76",  -- 118
        26742 => X"6D",  -- 109
        26743 => X"68",  -- 104
        26744 => X"60",  -- 96
        26745 => X"54",  -- 84
        26746 => X"43",  -- 67
        26747 => X"2C",  -- 44
        26748 => X"15",  -- 21
        26749 => X"0E",  -- 14
        26750 => X"1D",  -- 29
        26751 => X"34",  -- 52
        26752 => X"61",  -- 97
        26753 => X"6F",  -- 111
        26754 => X"78",  -- 120
        26755 => X"77",  -- 119
        26756 => X"89",  -- 137
        26757 => X"96",  -- 150
        26758 => X"90",  -- 144
        26759 => X"9E",  -- 158
        26760 => X"A6",  -- 166
        26761 => X"A6",  -- 166
        26762 => X"A8",  -- 168
        26763 => X"AD",  -- 173
        26764 => X"B6",  -- 182
        26765 => X"C0",  -- 192
        26766 => X"C4",  -- 196
        26767 => X"C3",  -- 195
        26768 => X"C0",  -- 192
        26769 => X"BF",  -- 191
        26770 => X"BE",  -- 190
        26771 => X"BE",  -- 190
        26772 => X"BF",  -- 191
        26773 => X"C0",  -- 192
        26774 => X"BE",  -- 190
        26775 => X"BB",  -- 187
        26776 => X"BE",  -- 190
        26777 => X"BD",  -- 189
        26778 => X"BD",  -- 189
        26779 => X"C2",  -- 194
        26780 => X"C8",  -- 200
        26781 => X"CB",  -- 203
        26782 => X"CA",  -- 202
        26783 => X"C7",  -- 199
        26784 => X"C4",  -- 196
        26785 => X"B2",  -- 178
        26786 => X"A2",  -- 162
        26787 => X"A4",  -- 164
        26788 => X"AD",  -- 173
        26789 => X"B4",  -- 180
        26790 => X"B7",  -- 183
        26791 => X"B9",  -- 185
        26792 => X"B5",  -- 181
        26793 => X"B8",  -- 184
        26794 => X"B9",  -- 185
        26795 => X"B4",  -- 180
        26796 => X"B0",  -- 176
        26797 => X"AC",  -- 172
        26798 => X"AA",  -- 170
        26799 => X"A6",  -- 166
        26800 => X"AB",  -- 171
        26801 => X"9C",  -- 156
        26802 => X"91",  -- 145
        26803 => X"92",  -- 146
        26804 => X"8F",  -- 143
        26805 => X"79",  -- 121
        26806 => X"53",  -- 83
        26807 => X"37",  -- 55
        26808 => X"3C",  -- 60
        26809 => X"3D",  -- 61
        26810 => X"47",  -- 71
        26811 => X"60",  -- 96
        26812 => X"7C",  -- 124
        26813 => X"93",  -- 147
        26814 => X"A0",  -- 160
        26815 => X"A7",  -- 167
        26816 => X"A8",  -- 168
        26817 => X"AE",  -- 174
        26818 => X"B0",  -- 176
        26819 => X"B9",  -- 185
        26820 => X"C7",  -- 199
        26821 => X"CC",  -- 204
        26822 => X"C9",  -- 201
        26823 => X"CC",  -- 204
        26824 => X"D1",  -- 209
        26825 => X"D1",  -- 209
        26826 => X"CD",  -- 205
        26827 => X"C9",  -- 201
        26828 => X"C4",  -- 196
        26829 => X"AE",  -- 174
        26830 => X"72",  -- 114
        26831 => X"34",  -- 52
        26832 => X"1D",  -- 29
        26833 => X"2C",  -- 44
        26834 => X"5B",  -- 91
        26835 => X"86",  -- 134
        26836 => X"90",  -- 144
        26837 => X"8E",  -- 142
        26838 => X"95",  -- 149
        26839 => X"99",  -- 153
        26840 => X"7B",  -- 123
        26841 => X"97",  -- 151
        26842 => X"A1",  -- 161
        26843 => X"92",  -- 146
        26844 => X"A6",  -- 166
        26845 => X"AB",  -- 171
        26846 => X"A8",  -- 168
        26847 => X"9F",  -- 159
        26848 => X"9B",  -- 155
        26849 => X"99",  -- 153
        26850 => X"9E",  -- 158
        26851 => X"A1",  -- 161
        26852 => X"9D",  -- 157
        26853 => X"A0",  -- 160
        26854 => X"A6",  -- 166
        26855 => X"A4",  -- 164
        26856 => X"AE",  -- 174
        26857 => X"9E",  -- 158
        26858 => X"90",  -- 144
        26859 => X"90",  -- 144
        26860 => X"9A",  -- 154
        26861 => X"A6",  -- 166
        26862 => X"A9",  -- 169
        26863 => X"AA",  -- 170
        26864 => X"AE",  -- 174
        26865 => X"A4",  -- 164
        26866 => X"A8",  -- 168
        26867 => X"BA",  -- 186
        26868 => X"C6",  -- 198
        26869 => X"C2",  -- 194
        26870 => X"BB",  -- 187
        26871 => X"B8",  -- 184
        26872 => X"C4",  -- 196
        26873 => X"C3",  -- 195
        26874 => X"BE",  -- 190
        26875 => X"B9",  -- 185
        26876 => X"AE",  -- 174
        26877 => X"A2",  -- 162
        26878 => X"97",  -- 151
        26879 => X"91",  -- 145
        26880 => X"69",  -- 105
        26881 => X"6A",  -- 106
        26882 => X"6B",  -- 107
        26883 => X"6D",  -- 109
        26884 => X"71",  -- 113
        26885 => X"71",  -- 113
        26886 => X"70",  -- 112
        26887 => X"6E",  -- 110
        26888 => X"68",  -- 104
        26889 => X"69",  -- 105
        26890 => X"69",  -- 105
        26891 => X"68",  -- 104
        26892 => X"68",  -- 104
        26893 => X"6B",  -- 107
        26894 => X"71",  -- 113
        26895 => X"78",  -- 120
        26896 => X"81",  -- 129
        26897 => X"8B",  -- 139
        26898 => X"96",  -- 150
        26899 => X"99",  -- 153
        26900 => X"9A",  -- 154
        26901 => X"99",  -- 153
        26902 => X"97",  -- 151
        26903 => X"93",  -- 147
        26904 => X"84",  -- 132
        26905 => X"7F",  -- 127
        26906 => X"79",  -- 121
        26907 => X"75",  -- 117
        26908 => X"6B",  -- 107
        26909 => X"60",  -- 96
        26910 => X"57",  -- 87
        26911 => X"55",  -- 85
        26912 => X"4C",  -- 76
        26913 => X"58",  -- 88
        26914 => X"50",  -- 80
        26915 => X"35",  -- 53
        26916 => X"35",  -- 53
        26917 => X"5E",  -- 94
        26918 => X"88",  -- 136
        26919 => X"9A",  -- 154
        26920 => X"85",  -- 133
        26921 => X"71",  -- 113
        26922 => X"51",  -- 81
        26923 => X"37",  -- 55
        26924 => X"26",  -- 38
        26925 => X"26",  -- 38
        26926 => X"3B",  -- 59
        26927 => X"50",  -- 80
        26928 => X"62",  -- 98
        26929 => X"67",  -- 103
        26930 => X"81",  -- 129
        26931 => X"94",  -- 148
        26932 => X"8E",  -- 142
        26933 => X"5D",  -- 93
        26934 => X"25",  -- 37
        26935 => X"1A",  -- 26
        26936 => X"04",  -- 4
        26937 => X"3A",  -- 58
        26938 => X"77",  -- 119
        26939 => X"98",  -- 152
        26940 => X"AB",  -- 171
        26941 => X"B7",  -- 183
        26942 => X"C7",  -- 199
        26943 => X"D3",  -- 211
        26944 => X"D5",  -- 213
        26945 => X"D0",  -- 208
        26946 => X"D1",  -- 209
        26947 => X"D4",  -- 212
        26948 => X"D3",  -- 211
        26949 => X"CC",  -- 204
        26950 => X"CF",  -- 207
        26951 => X"CF",  -- 207
        26952 => X"DF",  -- 223
        26953 => X"CC",  -- 204
        26954 => X"9E",  -- 158
        26955 => X"3A",  -- 58
        26956 => X"08",  -- 8
        26957 => X"0C",  -- 12
        26958 => X"02",  -- 2
        26959 => X"06",  -- 6
        26960 => X"0B",  -- 11
        26961 => X"2E",  -- 46
        26962 => X"70",  -- 112
        26963 => X"8E",  -- 142
        26964 => X"8D",  -- 141
        26965 => X"72",  -- 114
        26966 => X"4D",  -- 77
        26967 => X"1C",  -- 28
        26968 => X"10",  -- 16
        26969 => X"0C",  -- 12
        26970 => X"48",  -- 72
        26971 => X"57",  -- 87
        26972 => X"2B",  -- 43
        26973 => X"0B",  -- 11
        26974 => X"5E",  -- 94
        26975 => X"67",  -- 103
        26976 => X"60",  -- 96
        26977 => X"4E",  -- 78
        26978 => X"64",  -- 100
        26979 => X"83",  -- 131
        26980 => X"74",  -- 116
        26981 => X"70",  -- 112
        26982 => X"59",  -- 89
        26983 => X"57",  -- 87
        26984 => X"5A",  -- 90
        26985 => X"7F",  -- 127
        26986 => X"6E",  -- 110
        26987 => X"42",  -- 66
        26988 => X"1E",  -- 30
        26989 => X"0F",  -- 15
        26990 => X"13",  -- 19
        26991 => X"0B",  -- 11
        26992 => X"02",  -- 2
        26993 => X"09",  -- 9
        26994 => X"07",  -- 7
        26995 => X"15",  -- 21
        26996 => X"45",  -- 69
        26997 => X"B7",  -- 183
        26998 => X"E8",  -- 232
        26999 => X"D8",  -- 216
        27000 => X"E6",  -- 230
        27001 => X"E4",  -- 228
        27002 => X"E6",  -- 230
        27003 => X"E6",  -- 230
        27004 => X"E5",  -- 229
        27005 => X"E1",  -- 225
        27006 => X"DE",  -- 222
        27007 => X"DD",  -- 221
        27008 => X"E0",  -- 224
        27009 => X"C1",  -- 193
        27010 => X"BF",  -- 191
        27011 => X"C0",  -- 192
        27012 => X"A8",  -- 168
        27013 => X"96",  -- 150
        27014 => X"6A",  -- 106
        27015 => X"1E",  -- 30
        27016 => X"02",  -- 2
        27017 => X"0A",  -- 10
        27018 => X"25",  -- 37
        27019 => X"52",  -- 82
        27020 => X"81",  -- 129
        27021 => X"96",  -- 150
        27022 => X"96",  -- 150
        27023 => X"90",  -- 144
        27024 => X"8C",  -- 140
        27025 => X"79",  -- 121
        27026 => X"5E",  -- 94
        27027 => X"4D",  -- 77
        27028 => X"41",  -- 65
        27029 => X"34",  -- 52
        27030 => X"37",  -- 55
        27031 => X"4C",  -- 76
        27032 => X"5B",  -- 91
        27033 => X"92",  -- 146
        27034 => X"B0",  -- 176
        27035 => X"B5",  -- 181
        27036 => X"B0",  -- 176
        27037 => X"A2",  -- 162
        27038 => X"8A",  -- 138
        27039 => X"60",  -- 96
        27040 => X"61",  -- 97
        27041 => X"4F",  -- 79
        27042 => X"54",  -- 84
        27043 => X"8C",  -- 140
        27044 => X"B2",  -- 178
        27045 => X"B7",  -- 183
        27046 => X"B5",  -- 181
        27047 => X"A2",  -- 162
        27048 => X"6F",  -- 111
        27049 => X"5D",  -- 93
        27050 => X"59",  -- 89
        27051 => X"6A",  -- 106
        27052 => X"79",  -- 121
        27053 => X"7F",  -- 127
        27054 => X"7E",  -- 126
        27055 => X"7B",  -- 123
        27056 => X"6A",  -- 106
        27057 => X"70",  -- 112
        27058 => X"79",  -- 121
        27059 => X"7E",  -- 126
        27060 => X"7F",  -- 127
        27061 => X"79",  -- 121
        27062 => X"73",  -- 115
        27063 => X"6E",  -- 110
        27064 => X"67",  -- 103
        27065 => X"58",  -- 88
        27066 => X"42",  -- 66
        27067 => X"2C",  -- 44
        27068 => X"17",  -- 23
        27069 => X"0E",  -- 14
        27070 => X"1A",  -- 26
        27071 => X"2B",  -- 43
        27072 => X"40",  -- 64
        27073 => X"59",  -- 89
        27074 => X"6C",  -- 108
        27075 => X"6B",  -- 107
        27076 => X"81",  -- 129
        27077 => X"94",  -- 148
        27078 => X"86",  -- 134
        27079 => X"85",  -- 133
        27080 => X"99",  -- 153
        27081 => X"A5",  -- 165
        27082 => X"B0",  -- 176
        27083 => X"B1",  -- 177
        27084 => X"B0",  -- 176
        27085 => X"B9",  -- 185
        27086 => X"C7",  -- 199
        27087 => X"CF",  -- 207
        27088 => X"C8",  -- 200
        27089 => X"C4",  -- 196
        27090 => X"C1",  -- 193
        27091 => X"C0",  -- 192
        27092 => X"BF",  -- 191
        27093 => X"BE",  -- 190
        27094 => X"BD",  -- 189
        27095 => X"BD",  -- 189
        27096 => X"C2",  -- 194
        27097 => X"BF",  -- 191
        27098 => X"BD",  -- 189
        27099 => X"BC",  -- 188
        27100 => X"BE",  -- 190
        27101 => X"BD",  -- 189
        27102 => X"BA",  -- 186
        27103 => X"B7",  -- 183
        27104 => X"A8",  -- 168
        27105 => X"9C",  -- 156
        27106 => X"96",  -- 150
        27107 => X"A0",  -- 160
        27108 => X"A9",  -- 169
        27109 => X"AC",  -- 172
        27110 => X"AD",  -- 173
        27111 => X"B3",  -- 179
        27112 => X"BB",  -- 187
        27113 => X"BB",  -- 187
        27114 => X"B9",  -- 185
        27115 => X"B4",  -- 180
        27116 => X"B1",  -- 177
        27117 => X"B1",  -- 177
        27118 => X"AA",  -- 170
        27119 => X"A3",  -- 163
        27120 => X"A4",  -- 164
        27121 => X"A2",  -- 162
        27122 => X"A1",  -- 161
        27123 => X"9A",  -- 154
        27124 => X"88",  -- 136
        27125 => X"6B",  -- 107
        27126 => X"54",  -- 84
        27127 => X"47",  -- 71
        27128 => X"38",  -- 56
        27129 => X"3C",  -- 60
        27130 => X"40",  -- 64
        27131 => X"48",  -- 72
        27132 => X"63",  -- 99
        27133 => X"89",  -- 137
        27134 => X"A2",  -- 162
        27135 => X"A9",  -- 169
        27136 => X"AA",  -- 170
        27137 => X"B1",  -- 177
        27138 => X"B6",  -- 182
        27139 => X"BD",  -- 189
        27140 => X"CB",  -- 203
        27141 => X"CB",  -- 203
        27142 => X"C4",  -- 196
        27143 => X"C4",  -- 196
        27144 => X"CA",  -- 202
        27145 => X"CB",  -- 203
        27146 => X"C7",  -- 199
        27147 => X"C5",  -- 197
        27148 => X"BF",  -- 191
        27149 => X"9E",  -- 158
        27150 => X"5E",  -- 94
        27151 => X"2A",  -- 42
        27152 => X"20",  -- 32
        27153 => X"3B",  -- 59
        27154 => X"6B",  -- 107
        27155 => X"90",  -- 144
        27156 => X"90",  -- 144
        27157 => X"85",  -- 133
        27158 => X"8F",  -- 143
        27159 => X"A1",  -- 161
        27160 => X"96",  -- 150
        27161 => X"A1",  -- 161
        27162 => X"9C",  -- 156
        27163 => X"AA",  -- 170
        27164 => X"B4",  -- 180
        27165 => X"B1",  -- 177
        27166 => X"9D",  -- 157
        27167 => X"A4",  -- 164
        27168 => X"A6",  -- 166
        27169 => X"A0",  -- 160
        27170 => X"A1",  -- 161
        27171 => X"A2",  -- 162
        27172 => X"9E",  -- 158
        27173 => X"A2",  -- 162
        27174 => X"AA",  -- 170
        27175 => X"A9",  -- 169
        27176 => X"AC",  -- 172
        27177 => X"9A",  -- 154
        27178 => X"8D",  -- 141
        27179 => X"91",  -- 145
        27180 => X"9C",  -- 156
        27181 => X"A3",  -- 163
        27182 => X"A9",  -- 169
        27183 => X"AC",  -- 172
        27184 => X"AE",  -- 174
        27185 => X"A6",  -- 166
        27186 => X"A9",  -- 169
        27187 => X"BA",  -- 186
        27188 => X"C3",  -- 195
        27189 => X"BB",  -- 187
        27190 => X"B4",  -- 180
        27191 => X"B5",  -- 181
        27192 => X"B7",  -- 183
        27193 => X"BB",  -- 187
        27194 => X"BD",  -- 189
        27195 => X"BE",  -- 190
        27196 => X"BA",  -- 186
        27197 => X"B2",  -- 178
        27198 => X"AA",  -- 170
        27199 => X"A3",  -- 163
        27200 => X"66",  -- 102
        27201 => X"67",  -- 103
        27202 => X"69",  -- 105
        27203 => X"6E",  -- 110
        27204 => X"76",  -- 118
        27205 => X"7B",  -- 123
        27206 => X"7E",  -- 126
        27207 => X"7F",  -- 127
        27208 => X"78",  -- 120
        27209 => X"77",  -- 119
        27210 => X"75",  -- 117
        27211 => X"73",  -- 115
        27212 => X"70",  -- 112
        27213 => X"72",  -- 114
        27214 => X"75",  -- 117
        27215 => X"77",  -- 119
        27216 => X"7A",  -- 122
        27217 => X"81",  -- 129
        27218 => X"88",  -- 136
        27219 => X"8A",  -- 138
        27220 => X"8B",  -- 139
        27221 => X"8C",  -- 140
        27222 => X"89",  -- 137
        27223 => X"86",  -- 134
        27224 => X"78",  -- 120
        27225 => X"74",  -- 116
        27226 => X"73",  -- 115
        27227 => X"70",  -- 112
        27228 => X"6B",  -- 107
        27229 => X"63",  -- 99
        27230 => X"5F",  -- 95
        27231 => X"60",  -- 96
        27232 => X"68",  -- 104
        27233 => X"6B",  -- 107
        27234 => X"57",  -- 87
        27235 => X"3C",  -- 60
        27236 => X"4C",  -- 76
        27237 => X"7B",  -- 123
        27238 => X"8D",  -- 141
        27239 => X"82",  -- 130
        27240 => X"65",  -- 101
        27241 => X"4C",  -- 76
        27242 => X"31",  -- 49
        27243 => X"25",  -- 37
        27244 => X"20",  -- 32
        27245 => X"27",  -- 39
        27246 => X"3F",  -- 63
        27247 => X"57",  -- 87
        27248 => X"76",  -- 118
        27249 => X"75",  -- 117
        27250 => X"74",  -- 116
        27251 => X"5E",  -- 94
        27252 => X"3E",  -- 62
        27253 => X"26",  -- 38
        27254 => X"25",  -- 37
        27255 => X"48",  -- 72
        27256 => X"2C",  -- 44
        27257 => X"5E",  -- 94
        27258 => X"86",  -- 134
        27259 => X"9B",  -- 155
        27260 => X"AF",  -- 175
        27261 => X"BF",  -- 191
        27262 => X"C7",  -- 199
        27263 => X"CC",  -- 204
        27264 => X"CF",  -- 207
        27265 => X"D3",  -- 211
        27266 => X"D6",  -- 214
        27267 => X"D3",  -- 211
        27268 => X"D2",  -- 210
        27269 => X"CF",  -- 207
        27270 => X"DD",  -- 221
        27271 => X"CE",  -- 206
        27272 => X"CC",  -- 204
        27273 => X"78",  -- 120
        27274 => X"3B",  -- 59
        27275 => X"00",  -- 0
        27276 => X"05",  -- 5
        27277 => X"2A",  -- 42
        27278 => X"1F",  -- 31
        27279 => X"28",  -- 40
        27280 => X"42",  -- 66
        27281 => X"68",  -- 104
        27282 => X"80",  -- 128
        27283 => X"7B",  -- 123
        27284 => X"7F",  -- 127
        27285 => X"36",  -- 54
        27286 => X"0D",  -- 13
        27287 => X"11",  -- 17
        27288 => X"2B",  -- 43
        27289 => X"3F",  -- 63
        27290 => X"52",  -- 82
        27291 => X"4C",  -- 76
        27292 => X"0B",  -- 11
        27293 => X"1E",  -- 30
        27294 => X"6A",  -- 106
        27295 => X"78",  -- 120
        27296 => X"62",  -- 98
        27297 => X"2A",  -- 42
        27298 => X"22",  -- 34
        27299 => X"43",  -- 67
        27300 => X"61",  -- 97
        27301 => X"8E",  -- 142
        27302 => X"83",  -- 131
        27303 => X"85",  -- 133
        27304 => X"8B",  -- 139
        27305 => X"9D",  -- 157
        27306 => X"80",  -- 128
        27307 => X"6D",  -- 109
        27308 => X"5F",  -- 95
        27309 => X"41",  -- 65
        27310 => X"38",  -- 56
        27311 => X"2D",  -- 45
        27312 => X"1D",  -- 29
        27313 => X"13",  -- 19
        27314 => X"07",  -- 7
        27315 => X"05",  -- 5
        27316 => X"09",  -- 9
        27317 => X"61",  -- 97
        27318 => X"C1",  -- 193
        27319 => X"EF",  -- 239
        27320 => X"ED",  -- 237
        27321 => X"E8",  -- 232
        27322 => X"E3",  -- 227
        27323 => X"E6",  -- 230
        27324 => X"E8",  -- 232
        27325 => X"E8",  -- 232
        27326 => X"E1",  -- 225
        27327 => X"DB",  -- 219
        27328 => X"DE",  -- 222
        27329 => X"D1",  -- 209
        27330 => X"C9",  -- 201
        27331 => X"BB",  -- 187
        27332 => X"A8",  -- 168
        27333 => X"A1",  -- 161
        27334 => X"73",  -- 115
        27335 => X"27",  -- 39
        27336 => X"15",  -- 21
        27337 => X"15",  -- 21
        27338 => X"10",  -- 16
        27339 => X"18",  -- 24
        27340 => X"38",  -- 56
        27341 => X"5C",  -- 92
        27342 => X"7C",  -- 124
        27343 => X"97",  -- 151
        27344 => X"93",  -- 147
        27345 => X"7C",  -- 124
        27346 => X"61",  -- 97
        27347 => X"5A",  -- 90
        27348 => X"51",  -- 81
        27349 => X"39",  -- 57
        27350 => X"2F",  -- 47
        27351 => X"37",  -- 55
        27352 => X"40",  -- 64
        27353 => X"83",  -- 131
        27354 => X"B8",  -- 184
        27355 => X"CD",  -- 205
        27356 => X"C0",  -- 192
        27357 => X"9D",  -- 157
        27358 => X"8C",  -- 140
        27359 => X"85",  -- 133
        27360 => X"6C",  -- 108
        27361 => X"6C",  -- 108
        27362 => X"65",  -- 101
        27363 => X"83",  -- 131
        27364 => X"A9",  -- 169
        27365 => X"B3",  -- 179
        27366 => X"B5",  -- 181
        27367 => X"B1",  -- 177
        27368 => X"93",  -- 147
        27369 => X"79",  -- 121
        27370 => X"65",  -- 101
        27371 => X"67",  -- 103
        27372 => X"6A",  -- 106
        27373 => X"64",  -- 100
        27374 => X"5F",  -- 95
        27375 => X"63",  -- 99
        27376 => X"5D",  -- 93
        27377 => X"69",  -- 105
        27378 => X"79",  -- 121
        27379 => X"82",  -- 130
        27380 => X"84",  -- 132
        27381 => X"7E",  -- 126
        27382 => X"76",  -- 118
        27383 => X"72",  -- 114
        27384 => X"72",  -- 114
        27385 => X"60",  -- 96
        27386 => X"46",  -- 70
        27387 => X"30",  -- 48
        27388 => X"1B",  -- 27
        27389 => X"10",  -- 16
        27390 => X"16",  -- 22
        27391 => X"23",  -- 35
        27392 => X"28",  -- 40
        27393 => X"38",  -- 56
        27394 => X"45",  -- 69
        27395 => X"3E",  -- 62
        27396 => X"55",  -- 85
        27397 => X"76",  -- 118
        27398 => X"73",  -- 115
        27399 => X"6C",  -- 108
        27400 => X"7E",  -- 126
        27401 => X"96",  -- 150
        27402 => X"AE",  -- 174
        27403 => X"B3",  -- 179
        27404 => X"B2",  -- 178
        27405 => X"B9",  -- 185
        27406 => X"C6",  -- 198
        27407 => X"CE",  -- 206
        27408 => X"D5",  -- 213
        27409 => X"D0",  -- 208
        27410 => X"CD",  -- 205
        27411 => X"C9",  -- 201
        27412 => X"C3",  -- 195
        27413 => X"BE",  -- 190
        27414 => X"BD",  -- 189
        27415 => X"BF",  -- 191
        27416 => X"BF",  -- 191
        27417 => X"BF",  -- 191
        27418 => X"BD",  -- 189
        27419 => X"BB",  -- 187
        27420 => X"B8",  -- 184
        27421 => X"B7",  -- 183
        27422 => X"B5",  -- 181
        27423 => X"B2",  -- 178
        27424 => X"A0",  -- 160
        27425 => X"8D",  -- 141
        27426 => X"84",  -- 132
        27427 => X"96",  -- 150
        27428 => X"AC",  -- 172
        27429 => X"B7",  -- 183
        27430 => X"BA",  -- 186
        27431 => X"BD",  -- 189
        27432 => X"BA",  -- 186
        27433 => X"B8",  -- 184
        27434 => X"B6",  -- 182
        27435 => X"B4",  -- 180
        27436 => X"B7",  -- 183
        27437 => X"B8",  -- 184
        27438 => X"B5",  -- 181
        27439 => X"AE",  -- 174
        27440 => X"A1",  -- 161
        27441 => X"A8",  -- 168
        27442 => X"B0",  -- 176
        27443 => X"AB",  -- 171
        27444 => X"92",  -- 146
        27445 => X"6F",  -- 111
        27446 => X"4F",  -- 79
        27447 => X"41",  -- 65
        27448 => X"34",  -- 52
        27449 => X"2E",  -- 46
        27450 => X"2C",  -- 44
        27451 => X"3A",  -- 58
        27452 => X"53",  -- 83
        27453 => X"6E",  -- 110
        27454 => X"8B",  -- 139
        27455 => X"9F",  -- 159
        27456 => X"B1",  -- 177
        27457 => X"B9",  -- 185
        27458 => X"BC",  -- 188
        27459 => X"C4",  -- 196
        27460 => X"CD",  -- 205
        27461 => X"CC",  -- 204
        27462 => X"C5",  -- 197
        27463 => X"C4",  -- 196
        27464 => X"BF",  -- 191
        27465 => X"BF",  -- 191
        27466 => X"BC",  -- 188
        27467 => X"BD",  -- 189
        27468 => X"B6",  -- 182
        27469 => X"8D",  -- 141
        27470 => X"54",  -- 84
        27471 => X"34",  -- 52
        27472 => X"2E",  -- 46
        27473 => X"56",  -- 86
        27474 => X"81",  -- 129
        27475 => X"93",  -- 147
        27476 => X"99",  -- 153
        27477 => X"A2",  -- 162
        27478 => X"AB",  -- 171
        27479 => X"AF",  -- 175
        27480 => X"B0",  -- 176
        27481 => X"A8",  -- 168
        27482 => X"95",  -- 149
        27483 => X"B0",  -- 176
        27484 => X"B9",  -- 185
        27485 => X"B8",  -- 184
        27486 => X"A2",  -- 162
        27487 => X"B4",  -- 180
        27488 => X"AA",  -- 170
        27489 => X"A1",  -- 161
        27490 => X"A1",  -- 161
        27491 => X"A0",  -- 160
        27492 => X"9C",  -- 156
        27493 => X"A2",  -- 162
        27494 => X"AB",  -- 171
        27495 => X"AA",  -- 170
        27496 => X"A3",  -- 163
        27497 => X"93",  -- 147
        27498 => X"8A",  -- 138
        27499 => X"90",  -- 144
        27500 => X"9A",  -- 154
        27501 => X"9E",  -- 158
        27502 => X"A5",  -- 165
        27503 => X"AD",  -- 173
        27504 => X"B4",  -- 180
        27505 => X"B1",  -- 177
        27506 => X"B7",  -- 183
        27507 => X"C0",  -- 192
        27508 => X"C1",  -- 193
        27509 => X"B8",  -- 184
        27510 => X"B4",  -- 180
        27511 => X"B8",  -- 184
        27512 => X"B4",  -- 180
        27513 => X"B6",  -- 182
        27514 => X"B6",  -- 182
        27515 => X"B7",  -- 183
        27516 => X"B8",  -- 184
        27517 => X"B8",  -- 184
        27518 => X"B5",  -- 181
        27519 => X"AF",  -- 175
        27520 => X"69",  -- 105
        27521 => X"6A",  -- 106
        27522 => X"6D",  -- 109
        27523 => X"72",  -- 114
        27524 => X"79",  -- 121
        27525 => X"7E",  -- 126
        27526 => X"81",  -- 129
        27527 => X"82",  -- 130
        27528 => X"7F",  -- 127
        27529 => X"7B",  -- 123
        27530 => X"78",  -- 120
        27531 => X"74",  -- 116
        27532 => X"73",  -- 115
        27533 => X"72",  -- 114
        27534 => X"71",  -- 113
        27535 => X"71",  -- 113
        27536 => X"71",  -- 113
        27537 => X"74",  -- 116
        27538 => X"76",  -- 118
        27539 => X"75",  -- 117
        27540 => X"76",  -- 118
        27541 => X"78",  -- 120
        27542 => X"75",  -- 117
        27543 => X"71",  -- 113
        27544 => X"68",  -- 104
        27545 => X"67",  -- 103
        27546 => X"67",  -- 103
        27547 => X"68",  -- 104
        27548 => X"67",  -- 103
        27549 => X"65",  -- 101
        27550 => X"6A",  -- 106
        27551 => X"70",  -- 112
        27552 => X"7A",  -- 122
        27553 => X"6F",  -- 111
        27554 => X"53",  -- 83
        27555 => X"3E",  -- 62
        27556 => X"50",  -- 80
        27557 => X"73",  -- 115
        27558 => X"77",  -- 119
        27559 => X"61",  -- 97
        27560 => X"50",  -- 80
        27561 => X"3A",  -- 58
        27562 => X"2A",  -- 42
        27563 => X"2B",  -- 43
        27564 => X"34",  -- 52
        27565 => X"3F",  -- 63
        27566 => X"53",  -- 83
        27567 => X"68",  -- 104
        27568 => X"6C",  -- 108
        27569 => X"7C",  -- 124
        27570 => X"7C",  -- 124
        27571 => X"4C",  -- 76
        27572 => X"1E",  -- 30
        27573 => X"04",  -- 4
        27574 => X"01",  -- 1
        27575 => X"04",  -- 4
        27576 => X"37",  -- 55
        27577 => X"6D",  -- 109
        27578 => X"91",  -- 145
        27579 => X"9C",  -- 156
        27580 => X"B2",  -- 178
        27581 => X"C5",  -- 197
        27582 => X"C8",  -- 200
        27583 => X"C9",  -- 201
        27584 => X"C9",  -- 201
        27585 => X"D2",  -- 210
        27586 => X"D7",  -- 215
        27587 => X"D2",  -- 210
        27588 => X"D8",  -- 216
        27589 => X"D7",  -- 215
        27590 => X"D9",  -- 217
        27591 => X"A8",  -- 168
        27592 => X"7C",  -- 124
        27593 => X"2A",  -- 42
        27594 => X"06",  -- 6
        27595 => X"09",  -- 9
        27596 => X"22",  -- 34
        27597 => X"4C",  -- 76
        27598 => X"73",  -- 115
        27599 => X"98",  -- 152
        27600 => X"70",  -- 112
        27601 => X"51",  -- 81
        27602 => X"40",  -- 64
        27603 => X"47",  -- 71
        27604 => X"36",  -- 54
        27605 => X"06",  -- 6
        27606 => X"11",  -- 17
        27607 => X"58",  -- 88
        27608 => X"5A",  -- 90
        27609 => X"5B",  -- 91
        27610 => X"1E",  -- 30
        27611 => X"0E",  -- 14
        27612 => X"18",  -- 24
        27613 => X"4F",  -- 79
        27614 => X"64",  -- 100
        27615 => X"79",  -- 121
        27616 => X"68",  -- 104
        27617 => X"26",  -- 38
        27618 => X"06",  -- 6
        27619 => X"0A",  -- 10
        27620 => X"32",  -- 50
        27621 => X"77",  -- 119
        27622 => X"70",  -- 112
        27623 => X"72",  -- 114
        27624 => X"7E",  -- 126
        27625 => X"8D",  -- 141
        27626 => X"6E",  -- 110
        27627 => X"7F",  -- 127
        27628 => X"A3",  -- 163
        27629 => X"9C",  -- 156
        27630 => X"98",  -- 152
        27631 => X"87",  -- 135
        27632 => X"62",  -- 98
        27633 => X"31",  -- 49
        27634 => X"0D",  -- 13
        27635 => X"1D",  -- 29
        27636 => X"09",  -- 9
        27637 => X"0F",  -- 15
        27638 => X"54",  -- 84
        27639 => X"C0",  -- 192
        27640 => X"E5",  -- 229
        27641 => X"E4",  -- 228
        27642 => X"E3",  -- 227
        27643 => X"E4",  -- 228
        27644 => X"E7",  -- 231
        27645 => X"E9",  -- 233
        27646 => X"E4",  -- 228
        27647 => X"DF",  -- 223
        27648 => X"DA",  -- 218
        27649 => X"E4",  -- 228
        27650 => X"D2",  -- 210
        27651 => X"BC",  -- 188
        27652 => X"BD",  -- 189
        27653 => X"B6",  -- 182
        27654 => X"7B",  -- 123
        27655 => X"3C",  -- 60
        27656 => X"06",  -- 6
        27657 => X"0C",  -- 12
        27658 => X"08",  -- 8
        27659 => X"08",  -- 8
        27660 => X"15",  -- 21
        27661 => X"28",  -- 40
        27662 => X"53",  -- 83
        27663 => X"89",  -- 137
        27664 => X"A1",  -- 161
        27665 => X"91",  -- 145
        27666 => X"7D",  -- 125
        27667 => X"70",  -- 112
        27668 => X"67",  -- 103
        27669 => X"51",  -- 81
        27670 => X"42",  -- 66
        27671 => X"44",  -- 68
        27672 => X"53",  -- 83
        27673 => X"6C",  -- 108
        27674 => X"8B",  -- 139
        27675 => X"BB",  -- 187
        27676 => X"C5",  -- 197
        27677 => X"93",  -- 147
        27678 => X"74",  -- 116
        27679 => X"73",  -- 115
        27680 => X"6F",  -- 111
        27681 => X"71",  -- 113
        27682 => X"70",  -- 112
        27683 => X"8A",  -- 138
        27684 => X"A5",  -- 165
        27685 => X"AF",  -- 175
        27686 => X"B7",  -- 183
        27687 => X"B4",  -- 180
        27688 => X"A0",  -- 160
        27689 => X"87",  -- 135
        27690 => X"68",  -- 104
        27691 => X"5C",  -- 92
        27692 => X"60",  -- 96
        27693 => X"5E",  -- 94
        27694 => X"58",  -- 88
        27695 => X"59",  -- 89
        27696 => X"53",  -- 83
        27697 => X"64",  -- 100
        27698 => X"78",  -- 120
        27699 => X"85",  -- 133
        27700 => X"83",  -- 131
        27701 => X"7B",  -- 123
        27702 => X"72",  -- 114
        27703 => X"6F",  -- 111
        27704 => X"6C",  -- 108
        27705 => X"5A",  -- 90
        27706 => X"42",  -- 66
        27707 => X"2D",  -- 45
        27708 => X"1A",  -- 26
        27709 => X"0D",  -- 13
        27710 => X"13",  -- 19
        27711 => X"20",  -- 32
        27712 => X"24",  -- 36
        27713 => X"29",  -- 41
        27714 => X"34",  -- 52
        27715 => X"25",  -- 37
        27716 => X"25",  -- 37
        27717 => X"46",  -- 70
        27718 => X"56",  -- 86
        27719 => X"5A",  -- 90
        27720 => X"5B",  -- 91
        27721 => X"76",  -- 118
        27722 => X"90",  -- 144
        27723 => X"9C",  -- 156
        27724 => X"A1",  -- 161
        27725 => X"AD",  -- 173
        27726 => X"B5",  -- 181
        27727 => X"B8",  -- 184
        27728 => X"BB",  -- 187
        27729 => X"BC",  -- 188
        27730 => X"C0",  -- 192
        27731 => X"C1",  -- 193
        27732 => X"BE",  -- 190
        27733 => X"B9",  -- 185
        27734 => X"BC",  -- 188
        27735 => X"C2",  -- 194
        27736 => X"BC",  -- 188
        27737 => X"BE",  -- 190
        27738 => X"C2",  -- 194
        27739 => X"BF",  -- 191
        27740 => X"BB",  -- 187
        27741 => X"B8",  -- 184
        27742 => X"B7",  -- 183
        27743 => X"BA",  -- 186
        27744 => X"A1",  -- 161
        27745 => X"88",  -- 136
        27746 => X"7B",  -- 123
        27747 => X"8A",  -- 138
        27748 => X"A4",  -- 164
        27749 => X"B2",  -- 178
        27750 => X"B6",  -- 182
        27751 => X"BA",  -- 186
        27752 => X"BA",  -- 186
        27753 => X"BB",  -- 187
        27754 => X"BB",  -- 187
        27755 => X"BA",  -- 186
        27756 => X"BA",  -- 186
        27757 => X"BC",  -- 188
        27758 => X"BA",  -- 186
        27759 => X"B7",  -- 183
        27760 => X"B8",  -- 184
        27761 => X"B6",  -- 182
        27762 => X"B6",  -- 182
        27763 => X"B4",  -- 180
        27764 => X"A1",  -- 161
        27765 => X"73",  -- 115
        27766 => X"3B",  -- 59
        27767 => X"17",  -- 23
        27768 => X"25",  -- 37
        27769 => X"1D",  -- 29
        27770 => X"24",  -- 36
        27771 => X"3E",  -- 62
        27772 => X"5E",  -- 94
        27773 => X"7C",  -- 124
        27774 => X"9C",  -- 156
        27775 => X"B5",  -- 181
        27776 => X"B8",  -- 184
        27777 => X"BF",  -- 191
        27778 => X"C1",  -- 193
        27779 => X"C4",  -- 196
        27780 => X"CC",  -- 204
        27781 => X"CB",  -- 203
        27782 => X"C6",  -- 198
        27783 => X"C9",  -- 201
        27784 => X"CD",  -- 205
        27785 => X"C7",  -- 199
        27786 => X"BE",  -- 190
        27787 => X"B8",  -- 184
        27788 => X"A4",  -- 164
        27789 => X"6B",  -- 107
        27790 => X"35",  -- 53
        27791 => X"29",  -- 41
        27792 => X"40",  -- 64
        27793 => X"6F",  -- 111
        27794 => X"8F",  -- 143
        27795 => X"92",  -- 146
        27796 => X"9B",  -- 155
        27797 => X"AF",  -- 175
        27798 => X"B6",  -- 182
        27799 => X"B2",  -- 178
        27800 => X"B3",  -- 179
        27801 => X"A7",  -- 167
        27802 => X"95",  -- 149
        27803 => X"A1",  -- 161
        27804 => X"B7",  -- 183
        27805 => X"B8",  -- 184
        27806 => X"AE",  -- 174
        27807 => X"B8",  -- 184
        27808 => X"A9",  -- 169
        27809 => X"A1",  -- 161
        27810 => X"9E",  -- 158
        27811 => X"9D",  -- 157
        27812 => X"98",  -- 152
        27813 => X"9F",  -- 159
        27814 => X"A9",  -- 169
        27815 => X"A8",  -- 168
        27816 => X"9B",  -- 155
        27817 => X"8F",  -- 143
        27818 => X"8C",  -- 140
        27819 => X"94",  -- 148
        27820 => X"9B",  -- 155
        27821 => X"9C",  -- 156
        27822 => X"A4",  -- 164
        27823 => X"B1",  -- 177
        27824 => X"BA",  -- 186
        27825 => X"BE",  -- 190
        27826 => X"C2",  -- 194
        27827 => X"C2",  -- 194
        27828 => X"BA",  -- 186
        27829 => X"B0",  -- 176
        27830 => X"B2",  -- 178
        27831 => X"BA",  -- 186
        27832 => X"BB",  -- 187
        27833 => X"B9",  -- 185
        27834 => X"B5",  -- 181
        27835 => X"B2",  -- 178
        27836 => X"B2",  -- 178
        27837 => X"B4",  -- 180
        27838 => X"B1",  -- 177
        27839 => X"A9",  -- 169
        27840 => X"6A",  -- 106
        27841 => X"6B",  -- 107
        27842 => X"6D",  -- 109
        27843 => X"71",  -- 113
        27844 => X"75",  -- 117
        27845 => X"78",  -- 120
        27846 => X"78",  -- 120
        27847 => X"78",  -- 120
        27848 => X"7B",  -- 123
        27849 => X"77",  -- 119
        27850 => X"72",  -- 114
        27851 => X"6F",  -- 111
        27852 => X"6F",  -- 111
        27853 => X"6F",  -- 111
        27854 => X"6C",  -- 108
        27855 => X"6A",  -- 106
        27856 => X"6E",  -- 110
        27857 => X"6D",  -- 109
        27858 => X"6A",  -- 106
        27859 => X"67",  -- 103
        27860 => X"69",  -- 105
        27861 => X"6B",  -- 107
        27862 => X"68",  -- 104
        27863 => X"62",  -- 98
        27864 => X"62",  -- 98
        27865 => X"60",  -- 96
        27866 => X"61",  -- 97
        27867 => X"61",  -- 97
        27868 => X"63",  -- 99
        27869 => X"67",  -- 103
        27870 => X"71",  -- 113
        27871 => X"7C",  -- 124
        27872 => X"7D",  -- 125
        27873 => X"6E",  -- 110
        27874 => X"55",  -- 85
        27875 => X"48",  -- 72
        27876 => X"54",  -- 84
        27877 => X"6B",  -- 107
        27878 => X"6E",  -- 110
        27879 => X"62",  -- 98
        27880 => X"44",  -- 68
        27881 => X"32",  -- 50
        27882 => X"2C",  -- 44
        27883 => X"39",  -- 57
        27884 => X"4C",  -- 76
        27885 => X"59",  -- 89
        27886 => X"69",  -- 105
        27887 => X"7A",  -- 122
        27888 => X"74",  -- 116
        27889 => X"7B",  -- 123
        27890 => X"60",  -- 96
        27891 => X"21",  -- 33
        27892 => X"05",  -- 5
        27893 => X"0D",  -- 13
        27894 => X"0A",  -- 10
        27895 => X"09",  -- 9
        27896 => X"0F",  -- 15
        27897 => X"5B",  -- 91
        27898 => X"96",  -- 150
        27899 => X"AD",  -- 173
        27900 => X"C1",  -- 193
        27901 => X"CE",  -- 206
        27902 => X"CA",  -- 202
        27903 => X"C9",  -- 201
        27904 => X"CE",  -- 206
        27905 => X"D3",  -- 211
        27906 => X"D5",  -- 213
        27907 => X"CF",  -- 207
        27908 => X"DD",  -- 221
        27909 => X"D4",  -- 212
        27910 => X"BB",  -- 187
        27911 => X"65",  -- 101
        27912 => X"14",  -- 20
        27913 => X"02",  -- 2
        27914 => X"0C",  -- 12
        27915 => X"3E",  -- 62
        27916 => X"75",  -- 117
        27917 => X"AE",  -- 174
        27918 => X"CA",  -- 202
        27919 => X"AF",  -- 175
        27920 => X"4C",  -- 76
        27921 => X"0F",  -- 15
        27922 => X"16",  -- 22
        27923 => X"40",  -- 64
        27924 => X"0E",  -- 14
        27925 => X"0B",  -- 11
        27926 => X"3C",  -- 60
        27927 => X"6E",  -- 110
        27928 => X"72",  -- 114
        27929 => X"35",  -- 53
        27930 => X"06",  -- 6
        27931 => X"09",  -- 9
        27932 => X"40",  -- 64
        27933 => X"73",  -- 115
        27934 => X"78",  -- 120
        27935 => X"69",  -- 105
        27936 => X"76",  -- 118
        27937 => X"38",  -- 56
        27938 => X"0F",  -- 15
        27939 => X"07",  -- 7
        27940 => X"2D",  -- 45
        27941 => X"69",  -- 105
        27942 => X"41",  -- 65
        27943 => X"2A",  -- 42
        27944 => X"4B",  -- 75
        27945 => X"63",  -- 99
        27946 => X"3B",  -- 59
        27947 => X"3D",  -- 61
        27948 => X"6B",  -- 107
        27949 => X"92",  -- 146
        27950 => X"C0",  -- 192
        27951 => X"C9",  -- 201
        27952 => X"D0",  -- 208
        27953 => X"94",  -- 148
        27954 => X"52",  -- 82
        27955 => X"54",  -- 84
        27956 => X"3F",  -- 63
        27957 => X"14",  -- 20
        27958 => X"20",  -- 32
        27959 => X"7D",  -- 125
        27960 => X"DB",  -- 219
        27961 => X"E6",  -- 230
        27962 => X"EE",  -- 238
        27963 => X"EB",  -- 235
        27964 => X"E6",  -- 230
        27965 => X"E5",  -- 229
        27966 => X"E5",  -- 229
        27967 => X"E4",  -- 228
        27968 => X"E9",  -- 233
        27969 => X"D4",  -- 212
        27970 => X"DA",  -- 218
        27971 => X"D8",  -- 216
        27972 => X"BF",  -- 191
        27973 => X"B5",  -- 181
        27974 => X"8A",  -- 138
        27975 => X"35",  -- 53
        27976 => X"1C",  -- 28
        27977 => X"26",  -- 38
        27978 => X"25",  -- 37
        27979 => X"1E",  -- 30
        27980 => X"12",  -- 18
        27981 => X"0C",  -- 12
        27982 => X"35",  -- 53
        27983 => X"7A",  -- 122
        27984 => X"9B",  -- 155
        27985 => X"98",  -- 152
        27986 => X"87",  -- 135
        27987 => X"72",  -- 114
        27988 => X"66",  -- 102
        27989 => X"58",  -- 88
        27990 => X"4A",  -- 74
        27991 => X"4A",  -- 74
        27992 => X"5E",  -- 94
        27993 => X"79",  -- 121
        27994 => X"87",  -- 135
        27995 => X"A1",  -- 161
        27996 => X"A9",  -- 169
        27997 => X"8D",  -- 141
        27998 => X"7E",  -- 126
        27999 => X"81",  -- 129
        28000 => X"6C",  -- 108
        28001 => X"66",  -- 102
        28002 => X"6F",  -- 111
        28003 => X"91",  -- 145
        28004 => X"A6",  -- 166
        28005 => X"B3",  -- 179
        28006 => X"C2",  -- 194
        28007 => X"B5",  -- 181
        28008 => X"AD",  -- 173
        28009 => X"98",  -- 152
        28010 => X"71",  -- 113
        28011 => X"58",  -- 88
        28012 => X"58",  -- 88
        28013 => X"58",  -- 88
        28014 => X"4C",  -- 76
        28015 => X"40",  -- 64
        28016 => X"42",  -- 66
        28017 => X"56",  -- 86
        28018 => X"6F",  -- 111
        28019 => X"7E",  -- 126
        28020 => X"7C",  -- 124
        28021 => X"74",  -- 116
        28022 => X"6E",  -- 110
        28023 => X"6C",  -- 108
        28024 => X"59",  -- 89
        28025 => X"4B",  -- 75
        28026 => X"37",  -- 55
        28027 => X"26",  -- 38
        28028 => X"13",  -- 19
        28029 => X"0A",  -- 10
        28030 => X"12",  -- 18
        28031 => X"20",  -- 32
        28032 => X"1B",  -- 27
        28033 => X"27",  -- 39
        28034 => X"45",  -- 69
        28035 => X"37",  -- 55
        28036 => X"1D",  -- 29
        28037 => X"2B",  -- 43
        28038 => X"43",  -- 67
        28039 => X"54",  -- 84
        28040 => X"5D",  -- 93
        28041 => X"70",  -- 112
        28042 => X"87",  -- 135
        28043 => X"94",  -- 148
        28044 => X"A1",  -- 161
        28045 => X"B1",  -- 177
        28046 => X"B9",  -- 185
        28047 => X"B7",  -- 183
        28048 => X"C1",  -- 193
        28049 => X"C3",  -- 195
        28050 => X"C8",  -- 200
        28051 => X"C8",  -- 200
        28052 => X"BD",  -- 189
        28053 => X"B2",  -- 178
        28054 => X"B1",  -- 177
        28055 => X"B6",  -- 182
        28056 => X"C0",  -- 192
        28057 => X"C4",  -- 196
        28058 => X"C7",  -- 199
        28059 => X"C3",  -- 195
        28060 => X"BA",  -- 186
        28061 => X"B4",  -- 180
        28062 => X"B3",  -- 179
        28063 => X"B6",  -- 182
        28064 => X"AE",  -- 174
        28065 => X"99",  -- 153
        28066 => X"8D",  -- 141
        28067 => X"9B",  -- 155
        28068 => X"AD",  -- 173
        28069 => X"B7",  -- 183
        28070 => X"BF",  -- 191
        28071 => X"C8",  -- 200
        28072 => X"C9",  -- 201
        28073 => X"CD",  -- 205
        28074 => X"CD",  -- 205
        28075 => X"C4",  -- 196
        28076 => X"BC",  -- 188
        28077 => X"BA",  -- 186
        28078 => X"B7",  -- 183
        28079 => X"B6",  -- 182
        28080 => X"AF",  -- 175
        28081 => X"AA",  -- 170
        28082 => X"A7",  -- 167
        28083 => X"A6",  -- 166
        28084 => X"99",  -- 153
        28085 => X"75",  -- 117
        28086 => X"44",  -- 68
        28087 => X"24",  -- 36
        28088 => X"25",  -- 37
        28089 => X"20",  -- 32
        28090 => X"22",  -- 34
        28091 => X"32",  -- 50
        28092 => X"52",  -- 82
        28093 => X"77",  -- 119
        28094 => X"99",  -- 153
        28095 => X"AE",  -- 174
        28096 => X"C1",  -- 193
        28097 => X"C6",  -- 198
        28098 => X"C3",  -- 195
        28099 => X"C1",  -- 193
        28100 => X"C5",  -- 197
        28101 => X"C2",  -- 194
        28102 => X"BF",  -- 191
        28103 => X"C3",  -- 195
        28104 => X"C3",  -- 195
        28105 => X"BC",  -- 188
        28106 => X"B3",  -- 179
        28107 => X"AF",  -- 175
        28108 => X"99",  -- 153
        28109 => X"5C",  -- 92
        28110 => X"31",  -- 49
        28111 => X"32",  -- 50
        28112 => X"5C",  -- 92
        28113 => X"8C",  -- 140
        28114 => X"A8",  -- 168
        28115 => X"A6",  -- 166
        28116 => X"A7",  -- 167
        28117 => X"B2",  -- 178
        28118 => X"BA",  -- 186
        28119 => X"BE",  -- 190
        28120 => X"B9",  -- 185
        28121 => X"B1",  -- 177
        28122 => X"A5",  -- 165
        28123 => X"95",  -- 149
        28124 => X"B4",  -- 180
        28125 => X"B0",  -- 176
        28126 => X"AA",  -- 170
        28127 => X"A4",  -- 164
        28128 => X"AC",  -- 172
        28129 => X"A2",  -- 162
        28130 => X"9F",  -- 159
        28131 => X"9E",  -- 158
        28132 => X"99",  -- 153
        28133 => X"A0",  -- 160
        28134 => X"AA",  -- 170
        28135 => X"AA",  -- 170
        28136 => X"98",  -- 152
        28137 => X"8F",  -- 143
        28138 => X"8F",  -- 143
        28139 => X"99",  -- 153
        28140 => X"9F",  -- 159
        28141 => X"9D",  -- 157
        28142 => X"A8",  -- 168
        28143 => X"B9",  -- 185
        28144 => X"BE",  -- 190
        28145 => X"C3",  -- 195
        28146 => X"C6",  -- 198
        28147 => X"BF",  -- 191
        28148 => X"B1",  -- 177
        28149 => X"A9",  -- 169
        28150 => X"B1",  -- 177
        28151 => X"BB",  -- 187
        28152 => X"BC",  -- 188
        28153 => X"BB",  -- 187
        28154 => X"B6",  -- 182
        28155 => X"B3",  -- 179
        28156 => X"B3",  -- 179
        28157 => X"B4",  -- 180
        28158 => X"AD",  -- 173
        28159 => X"A2",  -- 162
        28160 => X"68",  -- 104
        28161 => X"67",  -- 103
        28162 => X"68",  -- 104
        28163 => X"6D",  -- 109
        28164 => X"72",  -- 114
        28165 => X"72",  -- 114
        28166 => X"6C",  -- 108
        28167 => X"66",  -- 102
        28168 => X"67",  -- 103
        28169 => X"69",  -- 105
        28170 => X"69",  -- 105
        28171 => X"68",  -- 104
        28172 => X"67",  -- 103
        28173 => X"6A",  -- 106
        28174 => X"72",  -- 114
        28175 => X"79",  -- 121
        28176 => X"7A",  -- 122
        28177 => X"79",  -- 121
        28178 => X"75",  -- 117
        28179 => X"70",  -- 112
        28180 => X"6D",  -- 109
        28181 => X"6B",  -- 107
        28182 => X"67",  -- 103
        28183 => X"64",  -- 100
        28184 => X"61",  -- 97
        28185 => X"62",  -- 98
        28186 => X"65",  -- 101
        28187 => X"65",  -- 101
        28188 => X"67",  -- 103
        28189 => X"6C",  -- 108
        28190 => X"75",  -- 117
        28191 => X"7D",  -- 125
        28192 => X"81",  -- 129
        28193 => X"72",  -- 114
        28194 => X"56",  -- 86
        28195 => X"47",  -- 71
        28196 => X"57",  -- 87
        28197 => X"70",  -- 112
        28198 => X"6E",  -- 110
        28199 => X"5C",  -- 92
        28200 => X"3C",  -- 60
        28201 => X"30",  -- 48
        28202 => X"37",  -- 55
        28203 => X"49",  -- 73
        28204 => X"54",  -- 84
        28205 => X"61",  -- 97
        28206 => X"73",  -- 115
        28207 => X"7C",  -- 124
        28208 => X"70",  -- 112
        28209 => X"73",  -- 115
        28210 => X"5F",  -- 95
        28211 => X"31",  -- 49
        28212 => X"1F",  -- 31
        28213 => X"14",  -- 20
        28214 => X"01",  -- 1
        28215 => X"02",  -- 2
        28216 => X"16",  -- 22
        28217 => X"59",  -- 89
        28218 => X"94",  -- 148
        28219 => X"A8",  -- 168
        28220 => X"BE",  -- 190
        28221 => X"CB",  -- 203
        28222 => X"C5",  -- 197
        28223 => X"CA",  -- 202
        28224 => X"D8",  -- 216
        28225 => X"C4",  -- 196
        28226 => X"C3",  -- 195
        28227 => X"DE",  -- 222
        28228 => X"D4",  -- 212
        28229 => X"CD",  -- 205
        28230 => X"76",  -- 118
        28231 => X"09",  -- 9
        28232 => X"0E",  -- 14
        28233 => X"4B",  -- 75
        28234 => X"59",  -- 89
        28235 => X"77",  -- 119
        28236 => X"D5",  -- 213
        28237 => X"D9",  -- 217
        28238 => X"D5",  -- 213
        28239 => X"8E",  -- 142
        28240 => X"23",  -- 35
        28241 => X"12",  -- 18
        28242 => X"66",  -- 102
        28243 => X"70",  -- 112
        28244 => X"18",  -- 24
        28245 => X"10",  -- 16
        28246 => X"1D",  -- 29
        28247 => X"68",  -- 104
        28248 => X"58",  -- 88
        28249 => X"27",  -- 39
        28250 => X"08",  -- 8
        28251 => X"2A",  -- 42
        28252 => X"67",  -- 103
        28253 => X"89",  -- 137
        28254 => X"6E",  -- 110
        28255 => X"6E",  -- 110
        28256 => X"77",  -- 119
        28257 => X"60",  -- 96
        28258 => X"26",  -- 38
        28259 => X"09",  -- 9
        28260 => X"30",  -- 48
        28261 => X"3A",  -- 58
        28262 => X"12",  -- 18
        28263 => X"0F",  -- 15
        28264 => X"12",  -- 18
        28265 => X"20",  -- 32
        28266 => X"13",  -- 19
        28267 => X"25",  -- 37
        28268 => X"16",  -- 22
        28269 => X"57",  -- 87
        28270 => X"BD",  -- 189
        28271 => X"D5",  -- 213
        28272 => X"DE",  -- 222
        28273 => X"C8",  -- 200
        28274 => X"C3",  -- 195
        28275 => X"B9",  -- 185
        28276 => X"A1",  -- 161
        28277 => X"6F",  -- 111
        28278 => X"17",  -- 23
        28279 => X"37",  -- 55
        28280 => X"C9",  -- 201
        28281 => X"D6",  -- 214
        28282 => X"F1",  -- 241
        28283 => X"E4",  -- 228
        28284 => X"E5",  -- 229
        28285 => X"DD",  -- 221
        28286 => X"E8",  -- 232
        28287 => X"DB",  -- 219
        28288 => X"DF",  -- 223
        28289 => X"E4",  -- 228
        28290 => X"DE",  -- 222
        28291 => X"DC",  -- 220
        28292 => X"C2",  -- 194
        28293 => X"AE",  -- 174
        28294 => X"95",  -- 149
        28295 => X"49",  -- 73
        28296 => X"22",  -- 34
        28297 => X"1D",  -- 29
        28298 => X"1A",  -- 26
        28299 => X"0F",  -- 15
        28300 => X"0C",  -- 12
        28301 => X"13",  -- 19
        28302 => X"23",  -- 35
        28303 => X"49",  -- 73
        28304 => X"89",  -- 137
        28305 => X"9F",  -- 159
        28306 => X"8D",  -- 141
        28307 => X"71",  -- 113
        28308 => X"63",  -- 99
        28309 => X"5E",  -- 94
        28310 => X"5C",  -- 92
        28311 => X"4E",  -- 78
        28312 => X"61",  -- 97
        28313 => X"64",  -- 100
        28314 => X"76",  -- 118
        28315 => X"9F",  -- 159
        28316 => X"B4",  -- 180
        28317 => X"9C",  -- 156
        28318 => X"81",  -- 129
        28319 => X"7C",  -- 124
        28320 => X"77",  -- 119
        28321 => X"6D",  -- 109
        28322 => X"71",  -- 113
        28323 => X"8D",  -- 141
        28324 => X"A9",  -- 169
        28325 => X"B3",  -- 179
        28326 => X"B4",  -- 180
        28327 => X"B2",  -- 178
        28328 => X"B4",  -- 180
        28329 => X"A5",  -- 165
        28330 => X"89",  -- 137
        28331 => X"6E",  -- 110
        28332 => X"5E",  -- 94
        28333 => X"58",  -- 88
        28334 => X"4F",  -- 79
        28335 => X"44",  -- 68
        28336 => X"4C",  -- 76
        28337 => X"56",  -- 86
        28338 => X"60",  -- 96
        28339 => X"63",  -- 99
        28340 => X"69",  -- 105
        28341 => X"6D",  -- 109
        28342 => X"6D",  -- 109
        28343 => X"69",  -- 105
        28344 => X"5A",  -- 90
        28345 => X"52",  -- 82
        28346 => X"38",  -- 56
        28347 => X"1D",  -- 29
        28348 => X"10",  -- 16
        28349 => X"0C",  -- 12
        28350 => X"11",  -- 17
        28351 => X"1E",  -- 30
        28352 => X"27",  -- 39
        28353 => X"2C",  -- 44
        28354 => X"39",  -- 57
        28355 => X"38",  -- 56
        28356 => X"24",  -- 36
        28357 => X"1B",  -- 27
        28358 => X"2A",  -- 42
        28359 => X"39",  -- 57
        28360 => X"4E",  -- 78
        28361 => X"68",  -- 104
        28362 => X"7C",  -- 124
        28363 => X"8F",  -- 143
        28364 => X"A1",  -- 161
        28365 => X"A2",  -- 162
        28366 => X"A7",  -- 167
        28367 => X"BC",  -- 188
        28368 => X"B8",  -- 184
        28369 => X"B8",  -- 184
        28370 => X"BA",  -- 186
        28371 => X"BE",  -- 190
        28372 => X"C1",  -- 193
        28373 => X"C2",  -- 194
        28374 => X"C1",  -- 193
        28375 => X"C0",  -- 192
        28376 => X"BE",  -- 190
        28377 => X"BD",  -- 189
        28378 => X"BD",  -- 189
        28379 => X"C1",  -- 193
        28380 => X"C6",  -- 198
        28381 => X"C3",  -- 195
        28382 => X"BC",  -- 188
        28383 => X"B6",  -- 182
        28384 => X"AF",  -- 175
        28385 => X"9D",  -- 157
        28386 => X"97",  -- 151
        28387 => X"9E",  -- 158
        28388 => X"AA",  -- 170
        28389 => X"BC",  -- 188
        28390 => X"C7",  -- 199
        28391 => X"C2",  -- 194
        28392 => X"BA",  -- 186
        28393 => X"B9",  -- 185
        28394 => X"BC",  -- 188
        28395 => X"BE",  -- 190
        28396 => X"BC",  -- 188
        28397 => X"B7",  -- 183
        28398 => X"BA",  -- 186
        28399 => X"C0",  -- 192
        28400 => X"B8",  -- 184
        28401 => X"B0",  -- 176
        28402 => X"AA",  -- 170
        28403 => X"AC",  -- 172
        28404 => X"A5",  -- 165
        28405 => X"86",  -- 134
        28406 => X"55",  -- 85
        28407 => X"30",  -- 48
        28408 => X"2C",  -- 44
        28409 => X"26",  -- 38
        28410 => X"21",  -- 33
        28411 => X"2F",  -- 47
        28412 => X"57",  -- 87
        28413 => X"8A",  -- 138
        28414 => X"AE",  -- 174
        28415 => X"BD",  -- 189
        28416 => X"BC",  -- 188
        28417 => X"BE",  -- 190
        28418 => X"C0",  -- 192
        28419 => X"C3",  -- 195
        28420 => X"C5",  -- 197
        28421 => X"C5",  -- 197
        28422 => X"C4",  -- 196
        28423 => X"C4",  -- 196
        28424 => X"C5",  -- 197
        28425 => X"AF",  -- 175
        28426 => X"B3",  -- 179
        28427 => X"A5",  -- 165
        28428 => X"7F",  -- 127
        28429 => X"4B",  -- 75
        28430 => X"2D",  -- 45
        28431 => X"4D",  -- 77
        28432 => X"85",  -- 133
        28433 => X"A6",  -- 166
        28434 => X"9F",  -- 159
        28435 => X"A4",  -- 164
        28436 => X"AD",  -- 173
        28437 => X"B7",  -- 183
        28438 => X"A8",  -- 168
        28439 => X"BD",  -- 189
        28440 => X"B2",  -- 178
        28441 => X"A9",  -- 169
        28442 => X"AB",  -- 171
        28443 => X"AF",  -- 175
        28444 => X"A8",  -- 168
        28445 => X"B7",  -- 183
        28446 => X"9C",  -- 156
        28447 => X"A5",  -- 165
        28448 => X"A8",  -- 168
        28449 => X"A9",  -- 169
        28450 => X"A6",  -- 166
        28451 => X"A3",  -- 163
        28452 => X"A6",  -- 166
        28453 => X"AB",  -- 171
        28454 => X"A5",  -- 165
        28455 => X"99",  -- 153
        28456 => X"94",  -- 148
        28457 => X"95",  -- 149
        28458 => X"99",  -- 153
        28459 => X"A1",  -- 161
        28460 => X"A4",  -- 164
        28461 => X"A4",  -- 164
        28462 => X"A9",  -- 169
        28463 => X"AD",  -- 173
        28464 => X"BA",  -- 186
        28465 => X"C1",  -- 193
        28466 => X"BF",  -- 191
        28467 => X"AF",  -- 175
        28468 => X"A2",  -- 162
        28469 => X"A5",  -- 165
        28470 => X"AD",  -- 173
        28471 => X"AF",  -- 175
        28472 => X"C0",  -- 192
        28473 => X"C3",  -- 195
        28474 => X"C2",  -- 194
        28475 => X"BC",  -- 188
        28476 => X"B8",  -- 184
        28477 => X"B6",  -- 182
        28478 => X"AE",  -- 174
        28479 => X"A4",  -- 164
        28480 => X"64",  -- 100
        28481 => X"64",  -- 100
        28482 => X"65",  -- 101
        28483 => X"69",  -- 105
        28484 => X"6D",  -- 109
        28485 => X"6E",  -- 110
        28486 => X"6C",  -- 108
        28487 => X"69",  -- 105
        28488 => X"6A",  -- 106
        28489 => X"6B",  -- 107
        28490 => X"69",  -- 105
        28491 => X"64",  -- 100
        28492 => X"62",  -- 98
        28493 => X"6A",  -- 106
        28494 => X"7A",  -- 122
        28495 => X"87",  -- 135
        28496 => X"88",  -- 136
        28497 => X"84",  -- 132
        28498 => X"7A",  -- 122
        28499 => X"73",  -- 115
        28500 => X"6E",  -- 110
        28501 => X"6A",  -- 106
        28502 => X"66",  -- 102
        28503 => X"62",  -- 98
        28504 => X"61",  -- 97
        28505 => X"62",  -- 98
        28506 => X"64",  -- 100
        28507 => X"65",  -- 101
        28508 => X"64",  -- 100
        28509 => X"6A",  -- 106
        28510 => X"72",  -- 114
        28511 => X"78",  -- 120
        28512 => X"84",  -- 132
        28513 => X"76",  -- 118
        28514 => X"63",  -- 99
        28515 => X"5C",  -- 92
        28516 => X"63",  -- 99
        28517 => X"6E",  -- 110
        28518 => X"6C",  -- 108
        28519 => X"63",  -- 99
        28520 => X"4C",  -- 76
        28521 => X"40",  -- 64
        28522 => X"44",  -- 68
        28523 => X"55",  -- 85
        28524 => X"5C",  -- 92
        28525 => X"65",  -- 101
        28526 => X"71",  -- 113
        28527 => X"79",  -- 121
        28528 => X"90",  -- 144
        28529 => X"5F",  -- 95
        28530 => X"28",  -- 40
        28531 => X"0E",  -- 14
        28532 => X"27",  -- 39
        28533 => X"36",  -- 54
        28534 => X"20",  -- 32
        28535 => X"18",  -- 24
        28536 => X"21",  -- 33
        28537 => X"5A",  -- 90
        28538 => X"92",  -- 146
        28539 => X"AE",  -- 174
        28540 => X"C1",  -- 193
        28541 => X"C1",  -- 193
        28542 => X"BC",  -- 188
        28543 => X"CC",  -- 204
        28544 => X"CB",  -- 203
        28545 => X"D8",  -- 216
        28546 => X"D0",  -- 208
        28547 => X"D1",  -- 209
        28548 => X"C5",  -- 197
        28549 => X"92",  -- 146
        28550 => X"45",  -- 69
        28551 => X"23",  -- 35
        28552 => X"73",  -- 115
        28553 => X"AA",  -- 170
        28554 => X"C3",  -- 195
        28555 => X"C6",  -- 198
        28556 => X"E4",  -- 228
        28557 => X"D9",  -- 217
        28558 => X"DA",  -- 218
        28559 => X"81",  -- 129
        28560 => X"1E",  -- 30
        28561 => X"3C",  -- 60
        28562 => X"92",  -- 146
        28563 => X"8B",  -- 139
        28564 => X"25",  -- 37
        28565 => X"15",  -- 21
        28566 => X"1D",  -- 29
        28567 => X"36",  -- 54
        28568 => X"3A",  -- 58
        28569 => X"0D",  -- 13
        28570 => X"15",  -- 21
        28571 => X"4E",  -- 78
        28572 => X"75",  -- 117
        28573 => X"80",  -- 128
        28574 => X"6E",  -- 110
        28575 => X"71",  -- 113
        28576 => X"74",  -- 116
        28577 => X"75",  -- 117
        28578 => X"4C",  -- 76
        28579 => X"1E",  -- 30
        28580 => X"17",  -- 23
        28581 => X"17",  -- 23
        28582 => X"05",  -- 5
        28583 => X"1D",  -- 29
        28584 => X"1F",  -- 31
        28585 => X"2B",  -- 43
        28586 => X"27",  -- 39
        28587 => X"43",  -- 67
        28588 => X"1A",  -- 26
        28589 => X"2C",  -- 44
        28590 => X"97",  -- 151
        28591 => X"D8",  -- 216
        28592 => X"DD",  -- 221
        28593 => X"DF",  -- 223
        28594 => X"E1",  -- 225
        28595 => X"D9",  -- 217
        28596 => X"DB",  -- 219
        28597 => X"C0",  -- 192
        28598 => X"65",  -- 101
        28599 => X"44",  -- 68
        28600 => X"75",  -- 117
        28601 => X"CD",  -- 205
        28602 => X"E7",  -- 231
        28603 => X"DA",  -- 218
        28604 => X"DF",  -- 223
        28605 => X"EE",  -- 238
        28606 => X"DF",  -- 223
        28607 => X"E5",  -- 229
        28608 => X"E1",  -- 225
        28609 => X"E5",  -- 229
        28610 => X"DD",  -- 221
        28611 => X"DA",  -- 218
        28612 => X"C1",  -- 193
        28613 => X"AA",  -- 170
        28614 => X"8E",  -- 142
        28615 => X"43",  -- 67
        28616 => X"11",  -- 17
        28617 => X"0B",  -- 11
        28618 => X"0E",  -- 14
        28619 => X"08",  -- 8
        28620 => X"0A",  -- 10
        28621 => X"0E",  -- 14
        28622 => X"18",  -- 24
        28623 => X"38",  -- 56
        28624 => X"89",  -- 137
        28625 => X"A5",  -- 165
        28626 => X"9D",  -- 157
        28627 => X"8A",  -- 138
        28628 => X"77",  -- 119
        28629 => X"5E",  -- 94
        28630 => X"56",  -- 86
        28631 => X"56",  -- 86
        28632 => X"5C",  -- 92
        28633 => X"63",  -- 99
        28634 => X"79",  -- 121
        28635 => X"9B",  -- 155
        28636 => X"B2",  -- 178
        28637 => X"A5",  -- 165
        28638 => X"8D",  -- 141
        28639 => X"82",  -- 130
        28640 => X"80",  -- 128
        28641 => X"77",  -- 119
        28642 => X"7B",  -- 123
        28643 => X"91",  -- 145
        28644 => X"A2",  -- 162
        28645 => X"A8",  -- 168
        28646 => X"B1",  -- 177
        28647 => X"BA",  -- 186
        28648 => X"AC",  -- 172
        28649 => X"A6",  -- 166
        28650 => X"99",  -- 153
        28651 => X"8B",  -- 139
        28652 => X"7A",  -- 122
        28653 => X"65",  -- 101
        28654 => X"4C",  -- 76
        28655 => X"39",  -- 57
        28656 => X"3C",  -- 60
        28657 => X"41",  -- 65
        28658 => X"47",  -- 71
        28659 => X"4C",  -- 76
        28660 => X"51",  -- 81
        28661 => X"55",  -- 85
        28662 => X"59",  -- 89
        28663 => X"5C",  -- 92
        28664 => X"49",  -- 73
        28665 => X"44",  -- 68
        28666 => X"2F",  -- 47
        28667 => X"1B",  -- 27
        28668 => X"13",  -- 19
        28669 => X"0E",  -- 14
        28670 => X"11",  -- 17
        28671 => X"1A",  -- 26
        28672 => X"33",  -- 51
        28673 => X"31",  -- 49
        28674 => X"2E",  -- 46
        28675 => X"23",  -- 35
        28676 => X"19",  -- 25
        28677 => X"1E",  -- 30
        28678 => X"22",  -- 34
        28679 => X"1D",  -- 29
        28680 => X"36",  -- 54
        28681 => X"60",  -- 96
        28682 => X"7D",  -- 125
        28683 => X"8C",  -- 140
        28684 => X"A1",  -- 161
        28685 => X"AC",  -- 172
        28686 => X"A8",  -- 168
        28687 => X"A8",  -- 168
        28688 => X"B3",  -- 179
        28689 => X"B6",  -- 182
        28690 => X"B9",  -- 185
        28691 => X"BB",  -- 187
        28692 => X"BA",  -- 186
        28693 => X"B9",  -- 185
        28694 => X"B8",  -- 184
        28695 => X"BA",  -- 186
        28696 => X"BA",  -- 186
        28697 => X"BB",  -- 187
        28698 => X"BD",  -- 189
        28699 => X"BD",  -- 189
        28700 => X"BE",  -- 190
        28701 => X"BC",  -- 188
        28702 => X"B7",  -- 183
        28703 => X"B3",  -- 179
        28704 => X"A8",  -- 168
        28705 => X"96",  -- 150
        28706 => X"93",  -- 147
        28707 => X"A1",  -- 161
        28708 => X"A6",  -- 166
        28709 => X"AC",  -- 172
        28710 => X"B6",  -- 182
        28711 => X"BC",  -- 188
        28712 => X"C1",  -- 193
        28713 => X"BD",  -- 189
        28714 => X"BF",  -- 191
        28715 => X"C4",  -- 196
        28716 => X"C5",  -- 197
        28717 => X"C4",  -- 196
        28718 => X"C6",  -- 198
        28719 => X"C8",  -- 200
        28720 => X"D2",  -- 210
        28721 => X"C9",  -- 201
        28722 => X"BF",  -- 191
        28723 => X"BA",  -- 186
        28724 => X"AF",  -- 175
        28725 => X"90",  -- 144
        28726 => X"5F",  -- 95
        28727 => X"36",  -- 54
        28728 => X"2B",  -- 43
        28729 => X"28",  -- 40
        28730 => X"2B",  -- 43
        28731 => X"3E",  -- 62
        28732 => X"62",  -- 98
        28733 => X"8B",  -- 139
        28734 => X"A8",  -- 168
        28735 => X"B7",  -- 183
        28736 => X"BC",  -- 188
        28737 => X"BD",  -- 189
        28738 => X"BF",  -- 191
        28739 => X"C2",  -- 194
        28740 => X"C4",  -- 196
        28741 => X"C4",  -- 196
        28742 => X"C6",  -- 198
        28743 => X"C5",  -- 197
        28744 => X"CD",  -- 205
        28745 => X"BC",  -- 188
        28746 => X"AA",  -- 170
        28747 => X"89",  -- 137
        28748 => X"64",  -- 100
        28749 => X"4B",  -- 75
        28750 => X"59",  -- 89
        28751 => X"8D",  -- 141
        28752 => X"98",  -- 152
        28753 => X"B1",  -- 177
        28754 => X"AD",  -- 173
        28755 => X"AA",  -- 170
        28756 => X"A2",  -- 162
        28757 => X"B8",  -- 184
        28758 => X"AF",  -- 175
        28759 => X"A6",  -- 166
        28760 => X"A6",  -- 166
        28761 => X"A6",  -- 166
        28762 => X"9F",  -- 159
        28763 => X"AB",  -- 171
        28764 => X"AF",  -- 175
        28765 => X"B4",  -- 180
        28766 => X"AD",  -- 173
        28767 => X"A4",  -- 164
        28768 => X"A8",  -- 168
        28769 => X"A9",  -- 169
        28770 => X"A8",  -- 168
        28771 => X"A9",  -- 169
        28772 => X"AC",  -- 172
        28773 => X"AB",  -- 171
        28774 => X"A3",  -- 163
        28775 => X"98",  -- 152
        28776 => X"92",  -- 146
        28777 => X"91",  -- 145
        28778 => X"97",  -- 151
        28779 => X"A0",  -- 160
        28780 => X"A7",  -- 167
        28781 => X"A8",  -- 168
        28782 => X"AA",  -- 170
        28783 => X"AC",  -- 172
        28784 => X"B4",  -- 180
        28785 => X"BE",  -- 190
        28786 => X"C1",  -- 193
        28787 => X"B3",  -- 179
        28788 => X"A7",  -- 167
        28789 => X"A6",  -- 166
        28790 => X"AB",  -- 171
        28791 => X"AE",  -- 174
        28792 => X"B4",  -- 180
        28793 => X"BD",  -- 189
        28794 => X"C1",  -- 193
        28795 => X"BE",  -- 190
        28796 => X"BE",  -- 190
        28797 => X"BE",  -- 190
        28798 => X"B7",  -- 183
        28799 => X"AC",  -- 172
        28800 => X"63",  -- 99
        28801 => X"64",  -- 100
        28802 => X"66",  -- 102
        28803 => X"67",  -- 103
        28804 => X"69",  -- 105
        28805 => X"6B",  -- 107
        28806 => X"6E",  -- 110
        28807 => X"71",  -- 113
        28808 => X"71",  -- 113
        28809 => X"70",  -- 112
        28810 => X"6C",  -- 108
        28811 => X"65",  -- 101
        28812 => X"62",  -- 98
        28813 => X"6B",  -- 107
        28814 => X"7F",  -- 127
        28815 => X"8F",  -- 143
        28816 => X"8B",  -- 139
        28817 => X"80",  -- 128
        28818 => X"73",  -- 115
        28819 => X"6A",  -- 106
        28820 => X"64",  -- 100
        28821 => X"60",  -- 96
        28822 => X"5D",  -- 93
        28823 => X"5B",  -- 91
        28824 => X"5A",  -- 90
        28825 => X"5B",  -- 91
        28826 => X"5D",  -- 93
        28827 => X"5B",  -- 91
        28828 => X"5D",  -- 93
        28829 => X"61",  -- 97
        28830 => X"6A",  -- 106
        28831 => X"6E",  -- 110
        28832 => X"70",  -- 112
        28833 => X"69",  -- 105
        28834 => X"5F",  -- 95
        28835 => X"5F",  -- 95
        28836 => X"6C",  -- 108
        28837 => X"77",  -- 119
        28838 => X"6C",  -- 108
        28839 => X"5B",  -- 91
        28840 => X"47",  -- 71
        28841 => X"3B",  -- 59
        28842 => X"43",  -- 67
        28843 => X"59",  -- 89
        28844 => X"64",  -- 100
        28845 => X"6C",  -- 108
        28846 => X"77",  -- 119
        28847 => X"7C",  -- 124
        28848 => X"74",  -- 116
        28849 => X"47",  -- 71
        28850 => X"1E",  -- 30
        28851 => X"08",  -- 8
        28852 => X"0B",  -- 11
        28853 => X"13",  -- 19
        28854 => X"1B",  -- 27
        28855 => X"38",  -- 56
        28856 => X"46",  -- 70
        28857 => X"78",  -- 120
        28858 => X"9D",  -- 157
        28859 => X"B0",  -- 176
        28860 => X"BC",  -- 188
        28861 => X"BB",  -- 187
        28862 => X"C2",  -- 194
        28863 => X"D6",  -- 214
        28864 => X"C7",  -- 199
        28865 => X"CC",  -- 204
        28866 => X"D8",  -- 216
        28867 => X"BF",  -- 191
        28868 => X"86",  -- 134
        28869 => X"5E",  -- 94
        28870 => X"7E",  -- 126
        28871 => X"AC",  -- 172
        28872 => X"BC",  -- 188
        28873 => X"D4",  -- 212
        28874 => X"E6",  -- 230
        28875 => X"E1",  -- 225
        28876 => X"E0",  -- 224
        28877 => X"D6",  -- 214
        28878 => X"CC",  -- 204
        28879 => X"53",  -- 83
        28880 => X"23",  -- 35
        28881 => X"7C",  -- 124
        28882 => X"9C",  -- 156
        28883 => X"6F",  -- 111
        28884 => X"30",  -- 48
        28885 => X"31",  -- 49
        28886 => X"39",  -- 57
        28887 => X"2F",  -- 47
        28888 => X"1A",  -- 26
        28889 => X"06",  -- 6
        28890 => X"31",  -- 49
        28891 => X"6F",  -- 111
        28892 => X"80",  -- 128
        28893 => X"79",  -- 121
        28894 => X"6E",  -- 110
        28895 => X"6A",  -- 106
        28896 => X"71",  -- 113
        28897 => X"89",  -- 137
        28898 => X"71",  -- 113
        28899 => X"3C",  -- 60
        28900 => X"09",  -- 9
        28901 => X"05",  -- 5
        28902 => X"06",  -- 6
        28903 => X"42",  -- 66
        28904 => X"55",  -- 85
        28905 => X"5F",  -- 95
        28906 => X"5C",  -- 92
        28907 => X"69",  -- 105
        28908 => X"34",  -- 52
        28909 => X"25",  -- 37
        28910 => X"8C",  -- 140
        28911 => X"DA",  -- 218
        28912 => X"D7",  -- 215
        28913 => X"DD",  -- 221
        28914 => X"DD",  -- 221
        28915 => X"D5",  -- 213
        28916 => X"E6",  -- 230
        28917 => X"DF",  -- 223
        28918 => X"AA",  -- 170
        28919 => X"69",  -- 105
        28920 => X"23",  -- 35
        28921 => X"65",  -- 101
        28922 => X"B6",  -- 182
        28923 => X"E2",  -- 226
        28924 => X"E4",  -- 228
        28925 => X"E4",  -- 228
        28926 => X"E4",  -- 228
        28927 => X"E1",  -- 225
        28928 => X"E9",  -- 233
        28929 => X"E9",  -- 233
        28930 => X"E0",  -- 224
        28931 => X"E2",  -- 226
        28932 => X"CC",  -- 204
        28933 => X"B4",  -- 180
        28934 => X"9A",  -- 154
        28935 => X"53",  -- 83
        28936 => X"0F",  -- 15
        28937 => X"07",  -- 7
        28938 => X"09",  -- 9
        28939 => X"07",  -- 7
        28940 => X"0B",  -- 11
        28941 => X"0B",  -- 11
        28942 => X"0F",  -- 15
        28943 => X"2B",  -- 43
        28944 => X"81",  -- 129
        28945 => X"AE",  -- 174
        28946 => X"AA",  -- 170
        28947 => X"98",  -- 152
        28948 => X"8A",  -- 138
        28949 => X"6B",  -- 107
        28950 => X"50",  -- 80
        28951 => X"45",  -- 69
        28952 => X"3F",  -- 63
        28953 => X"4D",  -- 77
        28954 => X"66",  -- 102
        28955 => X"87",  -- 135
        28956 => X"A6",  -- 166
        28957 => X"B3",  -- 179
        28958 => X"A9",  -- 169
        28959 => X"98",  -- 152
        28960 => X"86",  -- 134
        28961 => X"7E",  -- 126
        28962 => X"83",  -- 131
        28963 => X"96",  -- 150
        28964 => X"A0",  -- 160
        28965 => X"9F",  -- 159
        28966 => X"A9",  -- 169
        28967 => X"B9",  -- 185
        28968 => X"B0",  -- 176
        28969 => X"A4",  -- 164
        28970 => X"92",  -- 146
        28971 => X"85",  -- 133
        28972 => X"77",  -- 119
        28973 => X"68",  -- 104
        28974 => X"58",  -- 88
        28975 => X"4F",  -- 79
        28976 => X"3A",  -- 58
        28977 => X"33",  -- 51
        28978 => X"31",  -- 49
        28979 => X"35",  -- 53
        28980 => X"37",  -- 55
        28981 => X"38",  -- 56
        28982 => X"40",  -- 64
        28983 => X"4C",  -- 76
        28984 => X"44",  -- 68
        28985 => X"3E",  -- 62
        28986 => X"2C",  -- 44
        28987 => X"1A",  -- 26
        28988 => X"17",  -- 23
        28989 => X"15",  -- 21
        28990 => X"1B",  -- 27
        28991 => X"28",  -- 40
        28992 => X"45",  -- 69
        28993 => X"51",  -- 81
        28994 => X"47",  -- 71
        28995 => X"27",  -- 39
        28996 => X"15",  -- 21
        28997 => X"1E",  -- 30
        28998 => X"26",  -- 38
        28999 => X"24",  -- 36
        29000 => X"2E",  -- 46
        29001 => X"55",  -- 85
        29002 => X"77",  -- 119
        29003 => X"8F",  -- 143
        29004 => X"A9",  -- 169
        29005 => X"B6",  -- 182
        29006 => X"B1",  -- 177
        29007 => X"AD",  -- 173
        29008 => X"B2",  -- 178
        29009 => X"B7",  -- 183
        29010 => X"BB",  -- 187
        29011 => X"BA",  -- 186
        29012 => X"B6",  -- 182
        29013 => X"B3",  -- 179
        29014 => X"B4",  -- 180
        29015 => X"B6",  -- 182
        29016 => X"B1",  -- 177
        29017 => X"B4",  -- 180
        29018 => X"B8",  -- 184
        29019 => X"BA",  -- 186
        29020 => X"B9",  -- 185
        29021 => X"B7",  -- 183
        29022 => X"B6",  -- 182
        29023 => X"B5",  -- 181
        29024 => X"A5",  -- 165
        29025 => X"7F",  -- 127
        29026 => X"76",  -- 118
        29027 => X"93",  -- 147
        29028 => X"AD",  -- 173
        29029 => X"B5",  -- 181
        29030 => X"BA",  -- 186
        29031 => X"BA",  -- 186
        29032 => X"C6",  -- 198
        29033 => X"C2",  -- 194
        29034 => X"C0",  -- 192
        29035 => X"C6",  -- 198
        29036 => X"CA",  -- 202
        29037 => X"CB",  -- 203
        29038 => X"C9",  -- 201
        29039 => X"C8",  -- 200
        29040 => X"BF",  -- 191
        29041 => X"BE",  -- 190
        29042 => X"BD",  -- 189
        29043 => X"BD",  -- 189
        29044 => X"B3",  -- 179
        29045 => X"91",  -- 145
        29046 => X"56",  -- 86
        29047 => X"25",  -- 37
        29048 => X"28",  -- 40
        29049 => X"28",  -- 40
        29050 => X"30",  -- 48
        29051 => X"45",  -- 69
        29052 => X"66",  -- 102
        29053 => X"88",  -- 136
        29054 => X"A2",  -- 162
        29055 => X"B3",  -- 179
        29056 => X"BB",  -- 187
        29057 => X"BD",  -- 189
        29058 => X"C0",  -- 192
        29059 => X"C1",  -- 193
        29060 => X"C3",  -- 195
        29061 => X"C5",  -- 197
        29062 => X"C6",  -- 198
        29063 => X"C7",  -- 199
        29064 => X"C5",  -- 197
        29065 => X"BB",  -- 187
        29066 => X"96",  -- 150
        29067 => X"79",  -- 121
        29068 => X"63",  -- 99
        29069 => X"5F",  -- 95
        29070 => X"88",  -- 136
        29071 => X"B1",  -- 177
        29072 => X"AE",  -- 174
        29073 => X"B0",  -- 176
        29074 => X"B2",  -- 178
        29075 => X"B1",  -- 177
        29076 => X"A0",  -- 160
        29077 => X"B2",  -- 178
        29078 => X"B1",  -- 177
        29079 => X"9F",  -- 159
        29080 => X"A7",  -- 167
        29081 => X"AC",  -- 172
        29082 => X"9A",  -- 154
        29083 => X"A3",  -- 163
        29084 => X"B2",  -- 178
        29085 => X"AF",  -- 175
        29086 => X"BF",  -- 191
        29087 => X"AA",  -- 170
        29088 => X"A1",  -- 161
        29089 => X"A0",  -- 160
        29090 => X"A1",  -- 161
        29091 => X"A8",  -- 168
        29092 => X"A9",  -- 169
        29093 => X"A2",  -- 162
        29094 => X"97",  -- 151
        29095 => X"90",  -- 144
        29096 => X"92",  -- 146
        29097 => X"91",  -- 145
        29098 => X"95",  -- 149
        29099 => X"A1",  -- 161
        29100 => X"AA",  -- 170
        29101 => X"AA",  -- 170
        29102 => X"A9",  -- 169
        29103 => X"A9",  -- 169
        29104 => X"AF",  -- 175
        29105 => X"BB",  -- 187
        29106 => X"BD",  -- 189
        29107 => X"B1",  -- 177
        29108 => X"A4",  -- 164
        29109 => X"A4",  -- 164
        29110 => X"AB",  -- 171
        29111 => X"B0",  -- 176
        29112 => X"AE",  -- 174
        29113 => X"B7",  -- 183
        29114 => X"BE",  -- 190
        29115 => X"BF",  -- 191
        29116 => X"BF",  -- 191
        29117 => X"BE",  -- 190
        29118 => X"B5",  -- 181
        29119 => X"AA",  -- 170
        29120 => X"64",  -- 100
        29121 => X"67",  -- 103
        29122 => X"69",  -- 105
        29123 => X"67",  -- 103
        29124 => X"66",  -- 102
        29125 => X"68",  -- 104
        29126 => X"70",  -- 112
        29127 => X"76",  -- 118
        29128 => X"79",  -- 121
        29129 => X"76",  -- 118
        29130 => X"71",  -- 113
        29131 => X"6B",  -- 107
        29132 => X"69",  -- 105
        29133 => X"6E",  -- 110
        29134 => X"79",  -- 121
        29135 => X"83",  -- 131
        29136 => X"78",  -- 120
        29137 => X"6B",  -- 107
        29138 => X"5D",  -- 93
        29139 => X"57",  -- 87
        29140 => X"54",  -- 84
        29141 => X"54",  -- 84
        29142 => X"53",  -- 83
        29143 => X"53",  -- 83
        29144 => X"54",  -- 84
        29145 => X"57",  -- 87
        29146 => X"56",  -- 86
        29147 => X"55",  -- 85
        29148 => X"55",  -- 85
        29149 => X"5B",  -- 91
        29150 => X"61",  -- 97
        29151 => X"64",  -- 100
        29152 => X"5E",  -- 94
        29153 => X"5D",  -- 93
        29154 => X"56",  -- 86
        29155 => X"56",  -- 86
        29156 => X"6A",  -- 106
        29157 => X"76",  -- 118
        29158 => X"5B",  -- 91
        29159 => X"35",  -- 53
        29160 => X"32",  -- 50
        29161 => X"2C",  -- 44
        29162 => X"3C",  -- 60
        29163 => X"5A",  -- 90
        29164 => X"6B",  -- 107
        29165 => X"75",  -- 117
        29166 => X"81",  -- 129
        29167 => X"86",  -- 134
        29168 => X"68",  -- 104
        29169 => X"34",  -- 52
        29170 => X"13",  -- 19
        29171 => X"0B",  -- 11
        29172 => X"09",  -- 9
        29173 => X"01",  -- 1
        29174 => X"02",  -- 2
        29175 => X"22",  -- 34
        29176 => X"5D",  -- 93
        29177 => X"93",  -- 147
        29178 => X"AD",  -- 173
        29179 => X"B0",  -- 176
        29180 => X"B7",  -- 183
        29181 => X"BA",  -- 186
        29182 => X"C4",  -- 196
        29183 => X"CD",  -- 205
        29184 => X"D2",  -- 210
        29185 => X"D1",  -- 209
        29186 => X"C5",  -- 197
        29187 => X"77",  -- 119
        29188 => X"45",  -- 69
        29189 => X"5F",  -- 95
        29190 => X"BC",  -- 188
        29191 => X"E4",  -- 228
        29192 => X"C9",  -- 201
        29193 => X"CF",  -- 207
        29194 => X"D7",  -- 215
        29195 => X"DA",  -- 218
        29196 => X"DF",  -- 223
        29197 => X"DD",  -- 221
        29198 => X"CC",  -- 204
        29199 => X"5C",  -- 92
        29200 => X"4E",  -- 78
        29201 => X"A6",  -- 166
        29202 => X"7A",  -- 122
        29203 => X"44",  -- 68
        29204 => X"52",  -- 82
        29205 => X"67",  -- 103
        29206 => X"67",  -- 103
        29207 => X"4E",  -- 78
        29208 => X"12",  -- 18
        29209 => X"15",  -- 21
        29210 => X"4B",  -- 75
        29211 => X"71",  -- 113
        29212 => X"7C",  -- 124
        29213 => X"77",  -- 119
        29214 => X"6B",  -- 107
        29215 => X"5F",  -- 95
        29216 => X"71",  -- 113
        29217 => X"88",  -- 136
        29218 => X"7B",  -- 123
        29219 => X"57",  -- 87
        29220 => X"18",  -- 24
        29221 => X"08",  -- 8
        29222 => X"13",  -- 19
        29223 => X"5E",  -- 94
        29224 => X"7F",  -- 127
        29225 => X"92",  -- 146
        29226 => X"8B",  -- 139
        29227 => X"7B",  -- 123
        29228 => X"4D",  -- 77
        29229 => X"41",  -- 65
        29230 => X"A4",  -- 164
        29231 => X"DD",  -- 221
        29232 => X"DD",  -- 221
        29233 => X"D9",  -- 217
        29234 => X"D5",  -- 213
        29235 => X"CD",  -- 205
        29236 => X"D1",  -- 209
        29237 => X"C7",  -- 199
        29238 => X"D2",  -- 210
        29239 => X"AC",  -- 172
        29240 => X"54",  -- 84
        29241 => X"22",  -- 34
        29242 => X"5E",  -- 94
        29243 => X"A8",  -- 168
        29244 => X"E3",  -- 227
        29245 => X"CE",  -- 206
        29246 => X"E7",  -- 231
        29247 => X"E4",  -- 228
        29248 => X"E7",  -- 231
        29249 => X"E5",  -- 229
        29250 => X"DD",  -- 221
        29251 => X"E2",  -- 226
        29252 => X"D3",  -- 211
        29253 => X"C0",  -- 192
        29254 => X"AB",  -- 171
        29255 => X"65",  -- 101
        29256 => X"14",  -- 20
        29257 => X"08",  -- 8
        29258 => X"08",  -- 8
        29259 => X"07",  -- 7
        29260 => X"0B",  -- 11
        29261 => X"0C",  -- 12
        29262 => X"0E",  -- 14
        29263 => X"29",  -- 41
        29264 => X"7D",  -- 125
        29265 => X"B8",  -- 184
        29266 => X"B5",  -- 181
        29267 => X"99",  -- 153
        29268 => X"96",  -- 150
        29269 => X"86",  -- 134
        29270 => X"58",  -- 88
        29271 => X"2C",  -- 44
        29272 => X"20",  -- 32
        29273 => X"28",  -- 40
        29274 => X"3B",  -- 59
        29275 => X"58",  -- 88
        29276 => X"83",  -- 131
        29277 => X"AD",  -- 173
        29278 => X"B7",  -- 183
        29279 => X"A6",  -- 166
        29280 => X"8E",  -- 142
        29281 => X"85",  -- 133
        29282 => X"8A",  -- 138
        29283 => X"9F",  -- 159
        29284 => X"A8",  -- 168
        29285 => X"A3",  -- 163
        29286 => X"A6",  -- 166
        29287 => X"B3",  -- 179
        29288 => X"B7",  -- 183
        29289 => X"AC",  -- 172
        29290 => X"A3",  -- 163
        29291 => X"9D",  -- 157
        29292 => X"90",  -- 144
        29293 => X"7D",  -- 125
        29294 => X"6A",  -- 106
        29295 => X"5F",  -- 95
        29296 => X"4E",  -- 78
        29297 => X"3D",  -- 61
        29298 => X"33",  -- 51
        29299 => X"35",  -- 53
        29300 => X"30",  -- 48
        29301 => X"2A",  -- 42
        29302 => X"32",  -- 50
        29303 => X"42",  -- 66
        29304 => X"49",  -- 73
        29305 => X"43",  -- 67
        29306 => X"30",  -- 48
        29307 => X"1E",  -- 30
        29308 => X"18",  -- 24
        29309 => X"1B",  -- 27
        29310 => X"2B",  -- 43
        29311 => X"42",  -- 66
        29312 => X"46",  -- 70
        29313 => X"5E",  -- 94
        29314 => X"5C",  -- 92
        29315 => X"3D",  -- 61
        29316 => X"25",  -- 37
        29317 => X"22",  -- 34
        29318 => X"23",  -- 35
        29319 => X"23",  -- 35
        29320 => X"33",  -- 51
        29321 => X"44",  -- 68
        29322 => X"64",  -- 100
        29323 => X"8C",  -- 140
        29324 => X"A7",  -- 167
        29325 => X"B2",  -- 178
        29326 => X"B8",  -- 184
        29327 => X"C3",  -- 195
        29328 => X"BA",  -- 186
        29329 => X"BE",  -- 190
        29330 => X"C0",  -- 192
        29331 => X"BF",  -- 191
        29332 => X"BB",  -- 187
        29333 => X"B8",  -- 184
        29334 => X"B7",  -- 183
        29335 => X"B8",  -- 184
        29336 => X"B4",  -- 180
        29337 => X"B6",  -- 182
        29338 => X"B9",  -- 185
        29339 => X"BB",  -- 187
        29340 => X"BC",  -- 188
        29341 => X"B9",  -- 185
        29342 => X"B3",  -- 179
        29343 => X"AF",  -- 175
        29344 => X"9C",  -- 156
        29345 => X"75",  -- 117
        29346 => X"6B",  -- 107
        29347 => X"89",  -- 137
        29348 => X"AA",  -- 170
        29349 => X"BA",  -- 186
        29350 => X"C0",  -- 192
        29351 => X"C0",  -- 192
        29352 => X"C9",  -- 201
        29353 => X"C7",  -- 199
        29354 => X"C7",  -- 199
        29355 => X"C9",  -- 201
        29356 => X"CA",  -- 202
        29357 => X"C9",  -- 201
        29358 => X"C7",  -- 199
        29359 => X"C6",  -- 198
        29360 => X"B4",  -- 180
        29361 => X"B8",  -- 184
        29362 => X"BD",  -- 189
        29363 => X"C0",  -- 192
        29364 => X"BA",  -- 186
        29365 => X"9A",  -- 154
        29366 => X"63",  -- 99
        29367 => X"32",  -- 50
        29368 => X"2B",  -- 43
        29369 => X"27",  -- 39
        29370 => X"2C",  -- 44
        29371 => X"40",  -- 64
        29372 => X"60",  -- 96
        29373 => X"80",  -- 128
        29374 => X"A3",  -- 163
        29375 => X"BA",  -- 186
        29376 => X"BC",  -- 188
        29377 => X"BD",  -- 189
        29378 => X"BF",  -- 191
        29379 => X"C0",  -- 192
        29380 => X"C3",  -- 195
        29381 => X"C4",  -- 196
        29382 => X"C5",  -- 197
        29383 => X"C5",  -- 197
        29384 => X"C0",  -- 192
        29385 => X"AE",  -- 174
        29386 => X"7F",  -- 127
        29387 => X"79",  -- 121
        29388 => X"81",  -- 129
        29389 => X"85",  -- 133
        29390 => X"A2",  -- 162
        29391 => X"B2",  -- 178
        29392 => X"B7",  -- 183
        29393 => X"A9",  -- 169
        29394 => X"A8",  -- 168
        29395 => X"B1",  -- 177
        29396 => X"A9",  -- 169
        29397 => X"A6",  -- 166
        29398 => X"A8",  -- 168
        29399 => X"B1",  -- 177
        29400 => X"B1",  -- 177
        29401 => X"B0",  -- 176
        29402 => X"A3",  -- 163
        29403 => X"95",  -- 149
        29404 => X"A3",  -- 163
        29405 => X"A2",  -- 162
        29406 => X"B9",  -- 185
        29407 => X"AC",  -- 172
        29408 => X"9D",  -- 157
        29409 => X"97",  -- 151
        29410 => X"98",  -- 152
        29411 => X"A1",  -- 161
        29412 => X"A2",  -- 162
        29413 => X"97",  -- 151
        29414 => X"8E",  -- 142
        29415 => X"8A",  -- 138
        29416 => X"93",  -- 147
        29417 => X"94",  -- 148
        29418 => X"9B",  -- 155
        29419 => X"A4",  -- 164
        29420 => X"AB",  -- 171
        29421 => X"A9",  -- 169
        29422 => X"A9",  -- 169
        29423 => X"A8",  -- 168
        29424 => X"B2",  -- 178
        29425 => X"B9",  -- 185
        29426 => X"B6",  -- 182
        29427 => X"A8",  -- 168
        29428 => X"9D",  -- 157
        29429 => X"9E",  -- 158
        29430 => X"A9",  -- 169
        29431 => X"B3",  -- 179
        29432 => X"AE",  -- 174
        29433 => X"B5",  -- 181
        29434 => X"BA",  -- 186
        29435 => X"BA",  -- 186
        29436 => X"BB",  -- 187
        29437 => X"BC",  -- 188
        29438 => X"B4",  -- 180
        29439 => X"AB",  -- 171
        29440 => X"67",  -- 103
        29441 => X"6A",  -- 106
        29442 => X"6C",  -- 108
        29443 => X"69",  -- 105
        29444 => X"66",  -- 102
        29445 => X"68",  -- 104
        29446 => X"72",  -- 114
        29447 => X"7A",  -- 122
        29448 => X"7F",  -- 127
        29449 => X"7C",  -- 124
        29450 => X"78",  -- 120
        29451 => X"78",  -- 120
        29452 => X"7A",  -- 122
        29453 => X"7A",  -- 122
        29454 => X"77",  -- 119
        29455 => X"74",  -- 116
        29456 => X"64",  -- 100
        29457 => X"58",  -- 88
        29458 => X"4F",  -- 79
        29459 => X"4D",  -- 77
        29460 => X"50",  -- 80
        29461 => X"52",  -- 82
        29462 => X"54",  -- 84
        29463 => X"58",  -- 88
        29464 => X"61",  -- 97
        29465 => X"62",  -- 98
        29466 => X"60",  -- 96
        29467 => X"5B",  -- 91
        29468 => X"5B",  -- 91
        29469 => X"5F",  -- 95
        29470 => X"63",  -- 99
        29471 => X"62",  -- 98
        29472 => X"63",  -- 99
        29473 => X"5C",  -- 92
        29474 => X"59",  -- 89
        29475 => X"5E",  -- 94
        29476 => X"62",  -- 98
        29477 => X"53",  -- 83
        29478 => X"30",  -- 48
        29479 => X"13",  -- 19
        29480 => X"23",  -- 35
        29481 => X"24",  -- 36
        29482 => X"3C",  -- 60
        29483 => X"60",  -- 96
        29484 => X"73",  -- 115
        29485 => X"7C",  -- 124
        29486 => X"84",  -- 132
        29487 => X"87",  -- 135
        29488 => X"6C",  -- 108
        29489 => X"2C",  -- 44
        29490 => X"0C",  -- 12
        29491 => X"0F",  -- 15
        29492 => X"14",  -- 20
        29493 => X"09",  -- 9
        29494 => X"02",  -- 2
        29495 => X"17",  -- 23
        29496 => X"5E",  -- 94
        29497 => X"95",  -- 149
        29498 => X"AC",  -- 172
        29499 => X"B9",  -- 185
        29500 => X"C0",  -- 192
        29501 => X"B8",  -- 184
        29502 => X"BE",  -- 190
        29503 => X"C3",  -- 195
        29504 => X"CB",  -- 203
        29505 => X"C7",  -- 199
        29506 => X"8A",  -- 138
        29507 => X"3B",  -- 59
        29508 => X"68",  -- 104
        29509 => X"B0",  -- 176
        29510 => X"CE",  -- 206
        29511 => X"B8",  -- 184
        29512 => X"B5",  -- 181
        29513 => X"CE",  -- 206
        29514 => X"DA",  -- 218
        29515 => X"DD",  -- 221
        29516 => X"E2",  -- 226
        29517 => X"D9",  -- 217
        29518 => X"D4",  -- 212
        29519 => X"A1",  -- 161
        29520 => X"96",  -- 150
        29521 => X"94",  -- 148
        29522 => X"57",  -- 87
        29523 => X"57",  -- 87
        29524 => X"86",  -- 134
        29525 => X"90",  -- 144
        29526 => X"83",  -- 131
        29527 => X"57",  -- 87
        29528 => X"1A",  -- 26
        29529 => X"21",  -- 33
        29530 => X"44",  -- 68
        29531 => X"5F",  -- 95
        29532 => X"6E",  -- 110
        29533 => X"71",  -- 113
        29534 => X"63",  -- 99
        29535 => X"64",  -- 100
        29536 => X"74",  -- 116
        29537 => X"7C",  -- 124
        29538 => X"6E",  -- 110
        29539 => X"5F",  -- 95
        29540 => X"3E",  -- 62
        29541 => X"1D",  -- 29
        29542 => X"12",  -- 18
        29543 => X"4F",  -- 79
        29544 => X"74",  -- 116
        29545 => X"96",  -- 150
        29546 => X"A6",  -- 166
        29547 => X"88",  -- 136
        29548 => X"51",  -- 81
        29549 => X"3C",  -- 60
        29550 => X"AB",  -- 171
        29551 => X"DE",  -- 222
        29552 => X"DD",  -- 221
        29553 => X"D9",  -- 217
        29554 => X"D2",  -- 210
        29555 => X"C6",  -- 198
        29556 => X"B4",  -- 180
        29557 => X"A5",  -- 165
        29558 => X"D4",  -- 212
        29559 => X"CE",  -- 206
        29560 => X"B2",  -- 178
        29561 => X"64",  -- 100
        29562 => X"3E",  -- 62
        29563 => X"5B",  -- 91
        29564 => X"C4",  -- 196
        29565 => X"D8",  -- 216
        29566 => X"E1",  -- 225
        29567 => X"DD",  -- 221
        29568 => X"E4",  -- 228
        29569 => X"E3",  -- 227
        29570 => X"D8",  -- 216
        29571 => X"DD",  -- 221
        29572 => X"D0",  -- 208
        29573 => X"C3",  -- 195
        29574 => X"AF",  -- 175
        29575 => X"68",  -- 104
        29576 => X"0F",  -- 15
        29577 => X"03",  -- 3
        29578 => X"04",  -- 4
        29579 => X"06",  -- 6
        29580 => X"0A",  -- 10
        29581 => X"08",  -- 8
        29582 => X"0C",  -- 12
        29583 => X"29",  -- 41
        29584 => X"80",  -- 128
        29585 => X"BB",  -- 187
        29586 => X"BC",  -- 188
        29587 => X"A7",  -- 167
        29588 => X"A7",  -- 167
        29589 => X"99",  -- 153
        29590 => X"6D",  -- 109
        29591 => X"36",  -- 54
        29592 => X"18",  -- 24
        29593 => X"13",  -- 19
        29594 => X"18",  -- 24
        29595 => X"2A",  -- 42
        29596 => X"55",  -- 85
        29597 => X"8F",  -- 143
        29598 => X"AC",  -- 172
        29599 => X"A2",  -- 162
        29600 => X"A2",  -- 162
        29601 => X"94",  -- 148
        29602 => X"92",  -- 146
        29603 => X"A2",  -- 162
        29604 => X"AE",  -- 174
        29605 => X"AD",  -- 173
        29606 => X"AA",  -- 170
        29607 => X"AE",  -- 174
        29608 => X"B8",  -- 184
        29609 => X"AF",  -- 175
        29610 => X"A5",  -- 165
        29611 => X"9D",  -- 157
        29612 => X"8F",  -- 143
        29613 => X"7C",  -- 124
        29614 => X"69",  -- 105
        29615 => X"5E",  -- 94
        29616 => X"5D",  -- 93
        29617 => X"4A",  -- 74
        29618 => X"3C",  -- 60
        29619 => X"38",  -- 56
        29620 => X"31",  -- 49
        29621 => X"26",  -- 38
        29622 => X"2E",  -- 46
        29623 => X"3E",  -- 62
        29624 => X"43",  -- 67
        29625 => X"40",  -- 64
        29626 => X"30",  -- 48
        29627 => X"1E",  -- 30
        29628 => X"16",  -- 22
        29629 => X"19",  -- 25
        29630 => X"30",  -- 48
        29631 => X"4F",  -- 79
        29632 => X"53",  -- 83
        29633 => X"62",  -- 98
        29634 => X"61",  -- 97
        29635 => X"55",  -- 85
        29636 => X"4B",  -- 75
        29637 => X"37",  -- 55
        29638 => X"23",  -- 35
        29639 => X"1E",  -- 30
        29640 => X"2F",  -- 47
        29641 => X"36",  -- 54
        29642 => X"53",  -- 83
        29643 => X"78",  -- 120
        29644 => X"92",  -- 146
        29645 => X"A3",  -- 163
        29646 => X"B3",  -- 179
        29647 => X"C0",  -- 192
        29648 => X"C4",  -- 196
        29649 => X"C4",  -- 196
        29650 => X"C3",  -- 195
        29651 => X"C3",  -- 195
        29652 => X"C2",  -- 194
        29653 => X"C0",  -- 192
        29654 => X"BE",  -- 190
        29655 => X"BB",  -- 187
        29656 => X"C2",  -- 194
        29657 => X"BE",  -- 190
        29658 => X"BE",  -- 190
        29659 => X"C0",  -- 192
        29660 => X"C2",  -- 194
        29661 => X"BC",  -- 188
        29662 => X"B0",  -- 176
        29663 => X"A4",  -- 164
        29664 => X"92",  -- 146
        29665 => X"83",  -- 131
        29666 => X"86",  -- 134
        29667 => X"97",  -- 151
        29668 => X"A0",  -- 160
        29669 => X"AB",  -- 171
        29670 => X"B8",  -- 184
        29671 => X"C0",  -- 192
        29672 => X"C7",  -- 199
        29673 => X"CA",  -- 202
        29674 => X"CC",  -- 204
        29675 => X"CB",  -- 203
        29676 => X"CA",  -- 202
        29677 => X"C8",  -- 200
        29678 => X"C8",  -- 200
        29679 => X"C8",  -- 200
        29680 => X"C6",  -- 198
        29681 => X"C1",  -- 193
        29682 => X"BC",  -- 188
        29683 => X"B7",  -- 183
        29684 => X"AB",  -- 171
        29685 => X"91",  -- 145
        29686 => X"6B",  -- 107
        29687 => X"4C",  -- 76
        29688 => X"38",  -- 56
        29689 => X"2F",  -- 47
        29690 => X"2A",  -- 42
        29691 => X"36",  -- 54
        29692 => X"51",  -- 81
        29693 => X"7A",  -- 122
        29694 => X"A3",  -- 163
        29695 => X"C0",  -- 192
        29696 => X"BB",  -- 187
        29697 => X"BD",  -- 189
        29698 => X"BF",  -- 191
        29699 => X"C0",  -- 192
        29700 => X"C2",  -- 194
        29701 => X"C2",  -- 194
        29702 => X"C1",  -- 193
        29703 => X"C1",  -- 193
        29704 => X"BE",  -- 190
        29705 => X"A4",  -- 164
        29706 => X"74",  -- 116
        29707 => X"81",  -- 129
        29708 => X"9A",  -- 154
        29709 => X"9F",  -- 159
        29710 => X"B0",  -- 176
        29711 => X"B2",  -- 178
        29712 => X"AE",  -- 174
        29713 => X"B0",  -- 176
        29714 => X"A5",  -- 165
        29715 => X"A3",  -- 163
        29716 => X"AC",  -- 172
        29717 => X"9D",  -- 157
        29718 => X"9E",  -- 158
        29719 => X"BB",  -- 187
        29720 => X"B0",  -- 176
        29721 => X"A5",  -- 165
        29722 => X"AA",  -- 170
        29723 => X"8D",  -- 141
        29724 => X"93",  -- 147
        29725 => X"97",  -- 151
        29726 => X"9E",  -- 158
        29727 => X"A4",  -- 164
        29728 => X"A0",  -- 160
        29729 => X"98",  -- 152
        29730 => X"96",  -- 150
        29731 => X"9C",  -- 156
        29732 => X"9C",  -- 156
        29733 => X"95",  -- 149
        29734 => X"8F",  -- 143
        29735 => X"90",  -- 144
        29736 => X"92",  -- 146
        29737 => X"96",  -- 150
        29738 => X"A1",  -- 161
        29739 => X"AA",  -- 170
        29740 => X"AC",  -- 172
        29741 => X"AA",  -- 170
        29742 => X"AC",  -- 172
        29743 => X"B2",  -- 178
        29744 => X"B8",  -- 184
        29745 => X"BB",  -- 187
        29746 => X"B8",  -- 184
        29747 => X"AB",  -- 171
        29748 => X"9E",  -- 158
        29749 => X"9D",  -- 157
        29750 => X"A3",  -- 163
        29751 => X"A9",  -- 169
        29752 => X"AC",  -- 172
        29753 => X"B3",  -- 179
        29754 => X"B5",  -- 181
        29755 => X"B3",  -- 179
        29756 => X"B6",  -- 182
        29757 => X"BD",  -- 189
        29758 => X"BA",  -- 186
        29759 => X"B4",  -- 180
        29760 => X"6A",  -- 106
        29761 => X"6F",  -- 111
        29762 => X"71",  -- 113
        29763 => X"6F",  -- 111
        29764 => X"6C",  -- 108
        29765 => X"6F",  -- 111
        29766 => X"78",  -- 120
        29767 => X"81",  -- 129
        29768 => X"87",  -- 135
        29769 => X"83",  -- 131
        29770 => X"81",  -- 129
        29771 => X"84",  -- 132
        29772 => X"89",  -- 137
        29773 => X"86",  -- 134
        29774 => X"7B",  -- 123
        29775 => X"71",  -- 113
        29776 => X"5B",  -- 91
        29777 => X"55",  -- 85
        29778 => X"50",  -- 80
        29779 => X"55",  -- 85
        29780 => X"59",  -- 89
        29781 => X"5A",  -- 90
        29782 => X"60",  -- 96
        29783 => X"68",  -- 104
        29784 => X"74",  -- 116
        29785 => X"76",  -- 118
        29786 => X"71",  -- 113
        29787 => X"6A",  -- 106
        29788 => X"68",  -- 104
        29789 => X"6C",  -- 108
        29790 => X"6D",  -- 109
        29791 => X"68",  -- 104
        29792 => X"64",  -- 100
        29793 => X"59",  -- 89
        29794 => X"5C",  -- 92
        29795 => X"69",  -- 105
        29796 => X"52",  -- 82
        29797 => X"23",  -- 35
        29798 => X"0A",  -- 10
        29799 => X"0F",  -- 15
        29800 => X"12",  -- 18
        29801 => X"1A",  -- 26
        29802 => X"3E",  -- 62
        29803 => X"67",  -- 103
        29804 => X"79",  -- 121
        29805 => X"7F",  -- 127
        29806 => X"85",  -- 133
        29807 => X"89",  -- 137
        29808 => X"67",  -- 103
        29809 => X"2C",  -- 44
        29810 => X"13",  -- 19
        29811 => X"10",  -- 16
        29812 => X"09",  -- 9
        29813 => X"03",  -- 3
        29814 => X"0B",  -- 11
        29815 => X"28",  -- 40
        29816 => X"6A",  -- 106
        29817 => X"99",  -- 153
        29818 => X"A7",  -- 167
        29819 => X"BE",  -- 190
        29820 => X"C9",  -- 201
        29821 => X"BC",  -- 188
        29822 => X"C7",  -- 199
        29823 => X"D0",  -- 208
        29824 => X"B0",  -- 176
        29825 => X"6B",  -- 107
        29826 => X"4C",  -- 76
        29827 => X"6C",  -- 108
        29828 => X"B3",  -- 179
        29829 => X"DA",  -- 218
        29830 => X"D1",  -- 209
        29831 => X"A7",  -- 167
        29832 => X"A4",  -- 164
        29833 => X"CA",  -- 202
        29834 => X"D7",  -- 215
        29835 => X"DA",  -- 218
        29836 => X"E2",  -- 226
        29837 => X"DB",  -- 219
        29838 => X"DB",  -- 219
        29839 => X"CF",  -- 207
        29840 => X"BA",  -- 186
        29841 => X"59",  -- 89
        29842 => X"4D",  -- 77
        29843 => X"84",  -- 132
        29844 => X"9B",  -- 155
        29845 => X"94",  -- 148
        29846 => X"8A",  -- 138
        29847 => X"59",  -- 89
        29848 => X"22",  -- 34
        29849 => X"15",  -- 21
        29850 => X"28",  -- 40
        29851 => X"55",  -- 85
        29852 => X"58",  -- 88
        29853 => X"64",  -- 100
        29854 => X"60",  -- 96
        29855 => X"70",  -- 112
        29856 => X"78",  -- 120
        29857 => X"72",  -- 114
        29858 => X"5E",  -- 94
        29859 => X"4D",  -- 77
        29860 => X"57",  -- 87
        29861 => X"2C",  -- 44
        29862 => X"0B",  -- 11
        29863 => X"25",  -- 37
        29864 => X"63",  -- 99
        29865 => X"80",  -- 128
        29866 => X"B4",  -- 180
        29867 => X"A7",  -- 167
        29868 => X"58",  -- 88
        29869 => X"17",  -- 23
        29870 => X"95",  -- 149
        29871 => X"DE",  -- 222
        29872 => X"D9",  -- 217
        29873 => X"D8",  -- 216
        29874 => X"C7",  -- 199
        29875 => X"AD",  -- 173
        29876 => X"8F",  -- 143
        29877 => X"8D",  -- 141
        29878 => X"C1",  -- 193
        29879 => X"C9",  -- 201
        29880 => X"D6",  -- 214
        29881 => X"BA",  -- 186
        29882 => X"74",  -- 116
        29883 => X"4D",  -- 77
        29884 => X"58",  -- 88
        29885 => X"BD",  -- 189
        29886 => X"EA",  -- 234
        29887 => X"E5",  -- 229
        29888 => X"EA",  -- 234
        29889 => X"ED",  -- 237
        29890 => X"E1",  -- 225
        29891 => X"E0",  -- 224
        29892 => X"D4",  -- 212
        29893 => X"CB",  -- 203
        29894 => X"B2",  -- 178
        29895 => X"62",  -- 98
        29896 => X"11",  -- 17
        29897 => X"09",  -- 9
        29898 => X"0D",  -- 13
        29899 => X"0D",  -- 13
        29900 => X"0F",  -- 15
        29901 => X"0B",  -- 11
        29902 => X"11",  -- 17
        29903 => X"33",  -- 51
        29904 => X"8D",  -- 141
        29905 => X"B4",  -- 180
        29906 => X"BE",  -- 190
        29907 => X"BA",  -- 186
        29908 => X"AF",  -- 175
        29909 => X"9A",  -- 154
        29910 => X"80",  -- 128
        29911 => X"5B",  -- 91
        29912 => X"23",  -- 35
        29913 => X"10",  -- 16
        29914 => X"0B",  -- 11
        29915 => X"16",  -- 22
        29916 => X"35",  -- 53
        29917 => X"71",  -- 113
        29918 => X"A1",  -- 161
        29919 => X"A8",  -- 168
        29920 => X"B0",  -- 176
        29921 => X"A0",  -- 160
        29922 => X"95",  -- 149
        29923 => X"99",  -- 153
        29924 => X"A6",  -- 166
        29925 => X"AB",  -- 171
        29926 => X"AB",  -- 171
        29927 => X"AA",  -- 170
        29928 => X"CB",  -- 203
        29929 => X"C6",  -- 198
        29930 => X"BC",  -- 188
        29931 => X"AD",  -- 173
        29932 => X"A3",  -- 163
        29933 => X"9B",  -- 155
        29934 => X"91",  -- 145
        29935 => X"87",  -- 135
        29936 => X"5E",  -- 94
        29937 => X"4A",  -- 74
        29938 => X"39",  -- 57
        29939 => X"31",  -- 49
        29940 => X"27",  -- 39
        29941 => X"1E",  -- 30
        29942 => X"24",  -- 36
        29943 => X"34",  -- 52
        29944 => X"32",  -- 50
        29945 => X"2F",  -- 47
        29946 => X"24",  -- 36
        29947 => X"16",  -- 22
        29948 => X"11",  -- 17
        29949 => X"14",  -- 20
        29950 => X"2D",  -- 45
        29951 => X"4D",  -- 77
        29952 => X"6B",  -- 107
        29953 => X"72",  -- 114
        29954 => X"67",  -- 103
        29955 => X"59",  -- 89
        29956 => X"4E",  -- 78
        29957 => X"35",  -- 53
        29958 => X"29",  -- 41
        29959 => X"37",  -- 55
        29960 => X"26",  -- 38
        29961 => X"34",  -- 52
        29962 => X"4E",  -- 78
        29963 => X"66",  -- 102
        29964 => X"7B",  -- 123
        29965 => X"99",  -- 153
        29966 => X"AD",  -- 173
        29967 => X"AC",  -- 172
        29968 => X"C3",  -- 195
        29969 => X"C2",  -- 194
        29970 => X"C1",  -- 193
        29971 => X"C2",  -- 194
        29972 => X"C4",  -- 196
        29973 => X"C3",  -- 195
        29974 => X"C0",  -- 192
        29975 => X"BD",  -- 189
        29976 => X"C2",  -- 194
        29977 => X"BE",  -- 190
        29978 => X"BC",  -- 188
        29979 => X"C1",  -- 193
        29980 => X"C7",  -- 199
        29981 => X"C3",  -- 195
        29982 => X"B6",  -- 182
        29983 => X"AA",  -- 170
        29984 => X"98",  -- 152
        29985 => X"8C",  -- 140
        29986 => X"93",  -- 147
        29987 => X"A4",  -- 164
        29988 => X"AE",  -- 174
        29989 => X"B5",  -- 181
        29990 => X"BA",  -- 186
        29991 => X"B7",  -- 183
        29992 => X"C0",  -- 192
        29993 => X"C6",  -- 198
        29994 => X"CA",  -- 202
        29995 => X"C8",  -- 200
        29996 => X"C6",  -- 198
        29997 => X"C5",  -- 197
        29998 => X"C6",  -- 198
        29999 => X"C7",  -- 199
        30000 => X"C9",  -- 201
        30001 => X"C3",  -- 195
        30002 => X"BC",  -- 188
        30003 => X"B2",  -- 178
        30004 => X"99",  -- 153
        30005 => X"73",  -- 115
        30006 => X"52",  -- 82
        30007 => X"42",  -- 66
        30008 => X"3E",  -- 62
        30009 => X"35",  -- 53
        30010 => X"2A",  -- 42
        30011 => X"2B",  -- 43
        30012 => X"45",  -- 69
        30013 => X"72",  -- 114
        30014 => X"9F",  -- 159
        30015 => X"BA",  -- 186
        30016 => X"BB",  -- 187
        30017 => X"BD",  -- 189
        30018 => X"BF",  -- 191
        30019 => X"C0",  -- 192
        30020 => X"BF",  -- 191
        30021 => X"BF",  -- 191
        30022 => X"BD",  -- 189
        30023 => X"BC",  -- 188
        30024 => X"AB",  -- 171
        30025 => X"99",  -- 153
        30026 => X"82",  -- 130
        30027 => X"90",  -- 144
        30028 => X"A6",  -- 166
        30029 => X"A7",  -- 167
        30030 => X"A9",  -- 169
        30031 => X"AC",  -- 172
        30032 => X"A7",  -- 167
        30033 => X"BC",  -- 188
        30034 => X"AF",  -- 175
        30035 => X"95",  -- 149
        30036 => X"A5",  -- 165
        30037 => X"9D",  -- 157
        30038 => X"9C",  -- 156
        30039 => X"AE",  -- 174
        30040 => X"A8",  -- 168
        30041 => X"9E",  -- 158
        30042 => X"AD",  -- 173
        30043 => X"97",  -- 151
        30044 => X"91",  -- 145
        30045 => X"95",  -- 149
        30046 => X"8D",  -- 141
        30047 => X"9C",  -- 156
        30048 => X"A0",  -- 160
        30049 => X"99",  -- 153
        30050 => X"93",  -- 147
        30051 => X"94",  -- 148
        30052 => X"94",  -- 148
        30053 => X"94",  -- 148
        30054 => X"94",  -- 148
        30055 => X"97",  -- 151
        30056 => X"94",  -- 148
        30057 => X"9A",  -- 154
        30058 => X"A4",  -- 164
        30059 => X"AD",  -- 173
        30060 => X"AD",  -- 173
        30061 => X"AD",  -- 173
        30062 => X"B5",  -- 181
        30063 => X"BE",  -- 190
        30064 => X"BF",  -- 191
        30065 => X"C2",  -- 194
        30066 => X"C1",  -- 193
        30067 => X"B8",  -- 184
        30068 => X"AD",  -- 173
        30069 => X"A4",  -- 164
        30070 => X"A1",  -- 161
        30071 => X"A0",  -- 160
        30072 => X"AB",  -- 171
        30073 => X"B1",  -- 177
        30074 => X"B1",  -- 177
        30075 => X"AF",  -- 175
        30076 => X"B1",  -- 177
        30077 => X"B6",  -- 182
        30078 => X"B5",  -- 181
        30079 => X"AD",  -- 173
        30080 => X"64",  -- 100
        30081 => X"68",  -- 104
        30082 => X"6D",  -- 109
        30083 => X"6D",  -- 109
        30084 => X"6D",  -- 109
        30085 => X"70",  -- 112
        30086 => X"78",  -- 120
        30087 => X"7F",  -- 127
        30088 => X"83",  -- 131
        30089 => X"7E",  -- 126
        30090 => X"7A",  -- 122
        30091 => X"7C",  -- 124
        30092 => X"7F",  -- 127
        30093 => X"7C",  -- 124
        30094 => X"72",  -- 114
        30095 => X"6A",  -- 106
        30096 => X"58",  -- 88
        30097 => X"54",  -- 84
        30098 => X"57",  -- 87
        30099 => X"5D",  -- 93
        30100 => X"5D",  -- 93
        30101 => X"5B",  -- 91
        30102 => X"62",  -- 98
        30103 => X"6A",  -- 106
        30104 => X"71",  -- 113
        30105 => X"75",  -- 117
        30106 => X"71",  -- 113
        30107 => X"6A",  -- 106
        30108 => X"6A",  -- 106
        30109 => X"70",  -- 112
        30110 => X"71",  -- 113
        30111 => X"6B",  -- 107
        30112 => X"5F",  -- 95
        30113 => X"59",  -- 89
        30114 => X"60",  -- 96
        30115 => X"5F",  -- 95
        30116 => X"3E",  -- 62
        30117 => X"0F",  -- 15
        30118 => X"03",  -- 3
        30119 => X"13",  -- 19
        30120 => X"09",  -- 9
        30121 => X"18",  -- 24
        30122 => X"43",  -- 67
        30123 => X"6F",  -- 111
        30124 => X"80",  -- 128
        30125 => X"83",  -- 131
        30126 => X"89",  -- 137
        30127 => X"8E",  -- 142
        30128 => X"7D",  -- 125
        30129 => X"36",  -- 54
        30130 => X"13",  -- 19
        30131 => X"0C",  -- 12
        30132 => X"0B",  -- 11
        30133 => X"0F",  -- 15
        30134 => X"0E",  -- 14
        30135 => X"17",  -- 23
        30136 => X"68",  -- 104
        30137 => X"A7",  -- 167
        30138 => X"B1",  -- 177
        30139 => X"BB",  -- 187
        30140 => X"C5",  -- 197
        30141 => X"C3",  -- 195
        30142 => X"CB",  -- 203
        30143 => X"BA",  -- 186
        30144 => X"79",  -- 121
        30145 => X"1D",  -- 29
        30146 => X"44",  -- 68
        30147 => X"B9",  -- 185
        30148 => X"C3",  -- 195
        30149 => X"B1",  -- 177
        30150 => X"AE",  -- 174
        30151 => X"9F",  -- 159
        30152 => X"A9",  -- 169
        30153 => X"C9",  -- 201
        30154 => X"D7",  -- 215
        30155 => X"DC",  -- 220
        30156 => X"E2",  -- 226
        30157 => X"E7",  -- 231
        30158 => X"E3",  -- 227
        30159 => X"D0",  -- 208
        30160 => X"90",  -- 144
        30161 => X"41",  -- 65
        30162 => X"6E",  -- 110
        30163 => X"94",  -- 148
        30164 => X"95",  -- 149
        30165 => X"8E",  -- 142
        30166 => X"7F",  -- 127
        30167 => X"66",  -- 102
        30168 => X"20",  -- 32
        30169 => X"07",  -- 7
        30170 => X"1C",  -- 28
        30171 => X"57",  -- 87
        30172 => X"36",  -- 54
        30173 => X"5B",  -- 91
        30174 => X"65",  -- 101
        30175 => X"66",  -- 102
        30176 => X"76",  -- 118
        30177 => X"75",  -- 117
        30178 => X"52",  -- 82
        30179 => X"28",  -- 40
        30180 => X"52",  -- 82
        30181 => X"2F",  -- 47
        30182 => X"0B",  -- 11
        30183 => X"1B",  -- 27
        30184 => X"69",  -- 105
        30185 => X"61",  -- 97
        30186 => X"A7",  -- 167
        30187 => X"B8",  -- 184
        30188 => X"68",  -- 104
        30189 => X"09",  -- 9
        30190 => X"88",  -- 136
        30191 => X"DA",  -- 218
        30192 => X"DD",  -- 221
        30193 => X"DF",  -- 223
        30194 => X"C9",  -- 201
        30195 => X"AF",  -- 175
        30196 => X"87",  -- 135
        30197 => X"89",  -- 137
        30198 => X"AB",  -- 171
        30199 => X"C4",  -- 196
        30200 => X"DD",  -- 221
        30201 => X"DB",  -- 219
        30202 => X"B5",  -- 181
        30203 => X"78",  -- 120
        30204 => X"10",  -- 16
        30205 => X"5F",  -- 95
        30206 => X"B9",  -- 185
        30207 => X"DC",  -- 220
        30208 => X"E1",  -- 225
        30209 => X"EC",  -- 236
        30210 => X"E4",  -- 228
        30211 => X"E2",  -- 226
        30212 => X"D5",  -- 213
        30213 => X"D2",  -- 210
        30214 => X"B4",  -- 180
        30215 => X"5A",  -- 90
        30216 => X"19",  -- 25
        30217 => X"11",  -- 17
        30218 => X"14",  -- 20
        30219 => X"16",  -- 22
        30220 => X"18",  -- 24
        30221 => X"1F",  -- 31
        30222 => X"33",  -- 51
        30223 => X"63",  -- 99
        30224 => X"A0",  -- 160
        30225 => X"B4",  -- 180
        30226 => X"BD",  -- 189
        30227 => X"BD",  -- 189
        30228 => X"AA",  -- 170
        30229 => X"9E",  -- 158
        30230 => X"92",  -- 146
        30231 => X"6D",  -- 109
        30232 => X"2C",  -- 44
        30233 => X"12",  -- 18
        30234 => X"0D",  -- 13
        30235 => X"14",  -- 20
        30236 => X"20",  -- 32
        30237 => X"53",  -- 83
        30238 => X"93",  -- 147
        30239 => X"AA",  -- 170
        30240 => X"AA",  -- 170
        30241 => X"A6",  -- 166
        30242 => X"9D",  -- 157
        30243 => X"98",  -- 152
        30244 => X"9E",  -- 158
        30245 => X"A9",  -- 169
        30246 => X"AF",  -- 175
        30247 => X"AF",  -- 175
        30248 => X"AF",  -- 175
        30249 => X"BA",  -- 186
        30250 => X"C1",  -- 193
        30251 => X"BC",  -- 188
        30252 => X"B7",  -- 183
        30253 => X"B2",  -- 178
        30254 => X"A0",  -- 160
        30255 => X"8D",  -- 141
        30256 => X"69",  -- 105
        30257 => X"56",  -- 86
        30258 => X"3F",  -- 63
        30259 => X"2F",  -- 47
        30260 => X"21",  -- 33
        30261 => X"19",  -- 25
        30262 => X"1D",  -- 29
        30263 => X"29",  -- 41
        30264 => X"2D",  -- 45
        30265 => X"25",  -- 37
        30266 => X"15",  -- 21
        30267 => X"0C",  -- 12
        30268 => X"0F",  -- 15
        30269 => X"18",  -- 24
        30270 => X"34",  -- 52
        30271 => X"54",  -- 84
        30272 => X"72",  -- 114
        30273 => X"7A",  -- 122
        30274 => X"68",  -- 104
        30275 => X"50",  -- 80
        30276 => X"42",  -- 66
        30277 => X"2A",  -- 42
        30278 => X"20",  -- 32
        30279 => X"36",  -- 54
        30280 => X"26",  -- 38
        30281 => X"30",  -- 48
        30282 => X"4B",  -- 75
        30283 => X"63",  -- 99
        30284 => X"73",  -- 115
        30285 => X"91",  -- 145
        30286 => X"AA",  -- 170
        30287 => X"A9",  -- 169
        30288 => X"BA",  -- 186
        30289 => X"BC",  -- 188
        30290 => X"BE",  -- 190
        30291 => X"C0",  -- 192
        30292 => X"C0",  -- 192
        30293 => X"BF",  -- 191
        30294 => X"C0",  -- 192
        30295 => X"C0",  -- 192
        30296 => X"BC",  -- 188
        30297 => X"B9",  -- 185
        30298 => X"B8",  -- 184
        30299 => X"BC",  -- 188
        30300 => X"C3",  -- 195
        30301 => X"C3",  -- 195
        30302 => X"BB",  -- 187
        30303 => X"B3",  -- 179
        30304 => X"9E",  -- 158
        30305 => X"7F",  -- 127
        30306 => X"7D",  -- 125
        30307 => X"9D",  -- 157
        30308 => X"B8",  -- 184
        30309 => X"C2",  -- 194
        30310 => X"BE",  -- 190
        30311 => X"B7",  -- 183
        30312 => X"BE",  -- 190
        30313 => X"C3",  -- 195
        30314 => X"C6",  -- 198
        30315 => X"C5",  -- 197
        30316 => X"C4",  -- 196
        30317 => X"C5",  -- 197
        30318 => X"C3",  -- 195
        30319 => X"BF",  -- 191
        30320 => X"C5",  -- 197
        30321 => X"C1",  -- 193
        30322 => X"BF",  -- 191
        30323 => X"B8",  -- 184
        30324 => X"96",  -- 150
        30325 => X"62",  -- 98
        30326 => X"42",  -- 66
        30327 => X"3E",  -- 62
        30328 => X"3B",  -- 59
        30329 => X"39",  -- 57
        30330 => X"30",  -- 48
        30331 => X"2F",  -- 47
        30332 => X"49",  -- 73
        30333 => X"78",  -- 120
        30334 => X"9F",  -- 159
        30335 => X"B0",  -- 176
        30336 => X"BC",  -- 188
        30337 => X"BD",  -- 189
        30338 => X"C0",  -- 192
        30339 => X"C1",  -- 193
        30340 => X"BF",  -- 191
        30341 => X"BC",  -- 188
        30342 => X"B7",  -- 183
        30343 => X"B4",  -- 180
        30344 => X"A4",  -- 164
        30345 => X"9E",  -- 158
        30346 => X"9D",  -- 157
        30347 => X"9B",  -- 155
        30348 => X"A9",  -- 169
        30349 => X"AE",  -- 174
        30350 => X"A3",  -- 163
        30351 => X"A5",  -- 165
        30352 => X"A8",  -- 168
        30353 => X"B3",  -- 179
        30354 => X"B2",  -- 178
        30355 => X"9A",  -- 154
        30356 => X"A4",  -- 164
        30357 => X"9F",  -- 159
        30358 => X"A3",  -- 163
        30359 => X"A1",  -- 161
        30360 => X"A3",  -- 163
        30361 => X"A1",  -- 161
        30362 => X"A3",  -- 163
        30363 => X"A5",  -- 165
        30364 => X"99",  -- 153
        30365 => X"92",  -- 146
        30366 => X"8D",  -- 141
        30367 => X"97",  -- 151
        30368 => X"9B",  -- 155
        30369 => X"99",  -- 153
        30370 => X"91",  -- 145
        30371 => X"8B",  -- 139
        30372 => X"8C",  -- 140
        30373 => X"93",  -- 147
        30374 => X"99",  -- 153
        30375 => X"98",  -- 152
        30376 => X"9E",  -- 158
        30377 => X"A2",  -- 162
        30378 => X"A8",  -- 168
        30379 => X"AF",  -- 175
        30380 => X"B0",  -- 176
        30381 => X"B2",  -- 178
        30382 => X"B9",  -- 185
        30383 => X"C2",  -- 194
        30384 => X"BF",  -- 191
        30385 => X"C1",  -- 193
        30386 => X"C2",  -- 194
        30387 => X"C0",  -- 192
        30388 => X"BA",  -- 186
        30389 => X"B1",  -- 177
        30390 => X"AA",  -- 170
        30391 => X"A5",  -- 165
        30392 => X"AB",  -- 171
        30393 => X"B1",  -- 177
        30394 => X"B6",  -- 182
        30395 => X"B3",  -- 179
        30396 => X"B4",  -- 180
        30397 => X"B5",  -- 181
        30398 => X"AF",  -- 175
        30399 => X"A5",  -- 165
        30400 => X"55",  -- 85
        30401 => X"5B",  -- 91
        30402 => X"5F",  -- 95
        30403 => X"62",  -- 98
        30404 => X"63",  -- 99
        30405 => X"68",  -- 104
        30406 => X"6E",  -- 110
        30407 => X"75",  -- 117
        30408 => X"76",  -- 118
        30409 => X"70",  -- 112
        30410 => X"69",  -- 105
        30411 => X"65",  -- 101
        30412 => X"64",  -- 100
        30413 => X"62",  -- 98
        30414 => X"5E",  -- 94
        30415 => X"58",  -- 88
        30416 => X"56",  -- 86
        30417 => X"54",  -- 84
        30418 => X"56",  -- 86
        30419 => X"5E",  -- 94
        30420 => X"5C",  -- 92
        30421 => X"55",  -- 85
        30422 => X"59",  -- 89
        30423 => X"64",  -- 100
        30424 => X"62",  -- 98
        30425 => X"67",  -- 103
        30426 => X"65",  -- 101
        30427 => X"60",  -- 96
        30428 => X"63",  -- 99
        30429 => X"6C",  -- 108
        30430 => X"6E",  -- 110
        30431 => X"6A",  -- 106
        30432 => X"61",  -- 97
        30433 => X"69",  -- 105
        30434 => X"68",  -- 104
        30435 => X"50",  -- 80
        30436 => X"30",  -- 48
        30437 => X"18",  -- 24
        30438 => X"0E",  -- 14
        30439 => X"0E",  -- 14
        30440 => X"0F",  -- 15
        30441 => X"23",  -- 35
        30442 => X"51",  -- 81
        30443 => X"7E",  -- 126
        30444 => X"8A",  -- 138
        30445 => X"88",  -- 136
        30446 => X"8A",  -- 138
        30447 => X"8D",  -- 141
        30448 => X"8C",  -- 140
        30449 => X"50",  -- 80
        30450 => X"32",  -- 50
        30451 => X"23",  -- 35
        30452 => X"13",  -- 19
        30453 => X"0E",  -- 14
        30454 => X"09",  -- 9
        30455 => X"0B",  -- 11
        30456 => X"45",  -- 69
        30457 => X"AB",  -- 171
        30458 => X"C0",  -- 192
        30459 => X"B5",  -- 181
        30460 => X"BE",  -- 190
        30461 => X"C7",  -- 199
        30462 => X"BA",  -- 186
        30463 => X"7B",  -- 123
        30464 => X"2D",  -- 45
        30465 => X"21",  -- 33
        30466 => X"62",  -- 98
        30467 => X"CD",  -- 205
        30468 => X"C7",  -- 199
        30469 => X"AB",  -- 171
        30470 => X"9A",  -- 154
        30471 => X"A2",  -- 162
        30472 => X"AC",  -- 172
        30473 => X"C8",  -- 200
        30474 => X"E0",  -- 224
        30475 => X"DF",  -- 223
        30476 => X"D3",  -- 211
        30477 => X"DF",  -- 223
        30478 => X"DA",  -- 218
        30479 => X"BC",  -- 188
        30480 => X"4E",  -- 78
        30481 => X"55",  -- 85
        30482 => X"A2",  -- 162
        30483 => X"93",  -- 147
        30484 => X"96",  -- 150
        30485 => X"94",  -- 148
        30486 => X"6D",  -- 109
        30487 => X"6E",  -- 110
        30488 => X"1B",  -- 27
        30489 => X"07",  -- 7
        30490 => X"23",  -- 35
        30491 => X"5E",  -- 94
        30492 => X"1C",  -- 28
        30493 => X"5B",  -- 91
        30494 => X"6F",  -- 111
        30495 => X"52",  -- 82
        30496 => X"72",  -- 114
        30497 => X"79",  -- 121
        30498 => X"4D",  -- 77
        30499 => X"0A",  -- 10
        30500 => X"43",  -- 67
        30501 => X"30",  -- 48
        30502 => X"17",  -- 23
        30503 => X"28",  -- 40
        30504 => X"6B",  -- 107
        30505 => X"3F",  -- 63
        30506 => X"80",  -- 128
        30507 => X"AC",  -- 172
        30508 => X"73",  -- 115
        30509 => X"14",  -- 20
        30510 => X"91",  -- 145
        30511 => X"D4",  -- 212
        30512 => X"D3",  -- 211
        30513 => X"D6",  -- 214
        30514 => X"CD",  -- 205
        30515 => X"C4",  -- 196
        30516 => X"92",  -- 146
        30517 => X"85",  -- 133
        30518 => X"90",  -- 144
        30519 => X"BA",  -- 186
        30520 => X"CA",  -- 202
        30521 => X"D6",  -- 214
        30522 => X"DD",  -- 221
        30523 => X"C1",  -- 193
        30524 => X"56",  -- 86
        30525 => X"1F",  -- 31
        30526 => X"3F",  -- 63
        30527 => X"8D",  -- 141
        30528 => X"C9",  -- 201
        30529 => X"DC",  -- 220
        30530 => X"DA",  -- 218
        30531 => X"D7",  -- 215
        30532 => X"CE",  -- 206
        30533 => X"CF",  -- 207
        30534 => X"AF",  -- 175
        30535 => X"4D",  -- 77
        30536 => X"15",  -- 21
        30537 => X"0B",  -- 11
        30538 => X"10",  -- 16
        30539 => X"14",  -- 20
        30540 => X"21",  -- 33
        30541 => X"37",  -- 55
        30542 => X"61",  -- 97
        30543 => X"9F",  -- 159
        30544 => X"B5",  -- 181
        30545 => X"C0",  -- 192
        30546 => X"C0",  -- 192
        30547 => X"B6",  -- 182
        30548 => X"A6",  -- 166
        30549 => X"AE",  -- 174
        30550 => X"A5",  -- 165
        30551 => X"6A",  -- 106
        30552 => X"2F",  -- 47
        30553 => X"14",  -- 20
        30554 => X"0F",  -- 15
        30555 => X"12",  -- 18
        30556 => X"10",  -- 16
        30557 => X"36",  -- 54
        30558 => X"7A",  -- 122
        30559 => X"9E",  -- 158
        30560 => X"A1",  -- 161
        30561 => X"A8",  -- 168
        30562 => X"AA",  -- 170
        30563 => X"A2",  -- 162
        30564 => X"A3",  -- 163
        30565 => X"B0",  -- 176
        30566 => X"B9",  -- 185
        30567 => X"BA",  -- 186
        30568 => X"BB",  -- 187
        30569 => X"C3",  -- 195
        30570 => X"BF",  -- 191
        30571 => X"B1",  -- 177
        30572 => X"AD",  -- 173
        30573 => X"B3",  -- 179
        30574 => X"AF",  -- 175
        30575 => X"9F",  -- 159
        30576 => X"83",  -- 131
        30577 => X"70",  -- 112
        30578 => X"53",  -- 83
        30579 => X"3A",  -- 58
        30580 => X"26",  -- 38
        30581 => X"1B",  -- 27
        30582 => X"20",  -- 32
        30583 => X"28",  -- 40
        30584 => X"36",  -- 54
        30585 => X"27",  -- 39
        30586 => X"10",  -- 16
        30587 => X"08",  -- 8
        30588 => X"12",  -- 18
        30589 => X"22",  -- 34
        30590 => X"41",  -- 65
        30591 => X"64",  -- 100
        30592 => X"79",  -- 121
        30593 => X"7F",  -- 127
        30594 => X"6D",  -- 109
        30595 => X"5F",  -- 95
        30596 => X"60",  -- 96
        30597 => X"45",  -- 69
        30598 => X"20",  -- 32
        30599 => X"18",  -- 24
        30600 => X"2D",  -- 45
        30601 => X"27",  -- 39
        30602 => X"40",  -- 64
        30603 => X"65",  -- 101
        30604 => X"73",  -- 115
        30605 => X"87",  -- 135
        30606 => X"A6",  -- 166
        30607 => X"B7",  -- 183
        30608 => X"B2",  -- 178
        30609 => X"B7",  -- 183
        30610 => X"BD",  -- 189
        30611 => X"BF",  -- 191
        30612 => X"BC",  -- 188
        30613 => X"BB",  -- 187
        30614 => X"BE",  -- 190
        30615 => X"C2",  -- 194
        30616 => X"C1",  -- 193
        30617 => X"BE",  -- 190
        30618 => X"BC",  -- 188
        30619 => X"BA",  -- 186
        30620 => X"BA",  -- 186
        30621 => X"B9",  -- 185
        30622 => X"B4",  -- 180
        30623 => X"AF",  -- 175
        30624 => X"95",  -- 149
        30625 => X"70",  -- 112
        30626 => X"6B",  -- 107
        30627 => X"90",  -- 144
        30628 => X"AC",  -- 172
        30629 => X"B1",  -- 177
        30630 => X"B6",  -- 182
        30631 => X"BF",  -- 191
        30632 => X"C7",  -- 199
        30633 => X"C9",  -- 201
        30634 => X"C8",  -- 200
        30635 => X"C6",  -- 198
        30636 => X"C8",  -- 200
        30637 => X"CA",  -- 202
        30638 => X"C4",  -- 196
        30639 => X"BD",  -- 189
        30640 => X"C2",  -- 194
        30641 => X"BA",  -- 186
        30642 => X"B7",  -- 183
        30643 => X"AE",  -- 174
        30644 => X"89",  -- 137
        30645 => X"55",  -- 85
        30646 => X"42",  -- 66
        30647 => X"49",  -- 73
        30648 => X"39",  -- 57
        30649 => X"3E",  -- 62
        30650 => X"3B",  -- 59
        30651 => X"3B",  -- 59
        30652 => X"57",  -- 87
        30653 => X"88",  -- 136
        30654 => X"A9",  -- 169
        30655 => X"AF",  -- 175
        30656 => X"BB",  -- 187
        30657 => X"BD",  -- 189
        30658 => X"BF",  -- 191
        30659 => X"C0",  -- 192
        30660 => X"BF",  -- 191
        30661 => X"B9",  -- 185
        30662 => X"B4",  -- 180
        30663 => X"B1",  -- 177
        30664 => X"B7",  -- 183
        30665 => X"B2",  -- 178
        30666 => X"B0",  -- 176
        30667 => X"9A",  -- 154
        30668 => X"A3",  -- 163
        30669 => X"B9",  -- 185
        30670 => X"A9",  -- 169
        30671 => X"AA",  -- 170
        30672 => X"AD",  -- 173
        30673 => X"9F",  -- 159
        30674 => X"AC",  -- 172
        30675 => X"A9",  -- 169
        30676 => X"AB",  -- 171
        30677 => X"9F",  -- 159
        30678 => X"AA",  -- 170
        30679 => X"A0",  -- 160
        30680 => X"A2",  -- 162
        30681 => X"A6",  -- 166
        30682 => X"92",  -- 146
        30683 => X"A8",  -- 168
        30684 => X"97",  -- 151
        30685 => X"8B",  -- 139
        30686 => X"8F",  -- 143
        30687 => X"93",  -- 147
        30688 => X"9C",  -- 156
        30689 => X"9A",  -- 154
        30690 => X"93",  -- 147
        30691 => X"89",  -- 137
        30692 => X"8B",  -- 139
        30693 => X"96",  -- 150
        30694 => X"9D",  -- 157
        30695 => X"9C",  -- 156
        30696 => X"AB",  -- 171
        30697 => X"AA",  -- 170
        30698 => X"AB",  -- 171
        30699 => X"B0",  -- 176
        30700 => X"B3",  -- 179
        30701 => X"B3",  -- 179
        30702 => X"B9",  -- 185
        30703 => X"BE",  -- 190
        30704 => X"BD",  -- 189
        30705 => X"BC",  -- 188
        30706 => X"BD",  -- 189
        30707 => X"BE",  -- 190
        30708 => X"BD",  -- 189
        30709 => X"B8",  -- 184
        30710 => X"B4",  -- 180
        30711 => X"B2",  -- 178
        30712 => X"A7",  -- 167
        30713 => X"B1",  -- 177
        30714 => X"BA",  -- 186
        30715 => X"BD",  -- 189
        30716 => X"C1",  -- 193
        30717 => X"C1",  -- 193
        30718 => X"B7",  -- 183
        30719 => X"AC",  -- 172
        30720 => X"53",  -- 83
        30721 => X"52",  -- 82
        30722 => X"54",  -- 84
        30723 => X"55",  -- 85
        30724 => X"5A",  -- 90
        30725 => X"60",  -- 96
        30726 => X"65",  -- 101
        30727 => X"68",  -- 104
        30728 => X"67",  -- 103
        30729 => X"63",  -- 99
        30730 => X"5D",  -- 93
        30731 => X"56",  -- 86
        30732 => X"52",  -- 82
        30733 => X"4F",  -- 79
        30734 => X"4F",  -- 79
        30735 => X"50",  -- 80
        30736 => X"4F",  -- 79
        30737 => X"50",  -- 80
        30738 => X"50",  -- 80
        30739 => X"4F",  -- 79
        30740 => X"4F",  -- 79
        30741 => X"4C",  -- 76
        30742 => X"4A",  -- 74
        30743 => X"4A",  -- 74
        30744 => X"46",  -- 70
        30745 => X"47",  -- 71
        30746 => X"4B",  -- 75
        30747 => X"52",  -- 82
        30748 => X"5C",  -- 92
        30749 => X"62",  -- 98
        30750 => X"63",  -- 99
        30751 => X"61",  -- 97
        30752 => X"56",  -- 86
        30753 => X"67",  -- 103
        30754 => X"6E",  -- 110
        30755 => X"5A",  -- 90
        30756 => X"35",  -- 53
        30757 => X"17",  -- 23
        30758 => X"0B",  -- 11
        30759 => X"0B",  -- 11
        30760 => X"1A",  -- 26
        30761 => X"37",  -- 55
        30762 => X"68",  -- 104
        30763 => X"7E",  -- 126
        30764 => X"86",  -- 134
        30765 => X"8E",  -- 142
        30766 => X"8B",  -- 139
        30767 => X"86",  -- 134
        30768 => X"87",  -- 135
        30769 => X"73",  -- 115
        30770 => X"67",  -- 103
        30771 => X"61",  -- 97
        30772 => X"40",  -- 64
        30773 => X"15",  -- 21
        30774 => X"09",  -- 9
        30775 => X"17",  -- 23
        30776 => X"4E",  -- 78
        30777 => X"95",  -- 149
        30778 => X"BF",  -- 191
        30779 => X"C9",  -- 201
        30780 => X"A1",  -- 161
        30781 => X"83",  -- 131
        30782 => X"85",  -- 133
        30783 => X"5C",  -- 92
        30784 => X"11",  -- 17
        30785 => X"30",  -- 48
        30786 => X"8B",  -- 139
        30787 => X"C1",  -- 193
        30788 => X"C9",  -- 201
        30789 => X"A3",  -- 163
        30790 => X"73",  -- 115
        30791 => X"8C",  -- 140
        30792 => X"AD",  -- 173
        30793 => X"CE",  -- 206
        30794 => X"D6",  -- 214
        30795 => X"DD",  -- 221
        30796 => X"DE",  -- 222
        30797 => X"DF",  -- 223
        30798 => X"C9",  -- 201
        30799 => X"80",  -- 128
        30800 => X"28",  -- 40
        30801 => X"7B",  -- 123
        30802 => X"9F",  -- 159
        30803 => X"83",  -- 131
        30804 => X"65",  -- 101
        30805 => X"5A",  -- 90
        30806 => X"82",  -- 130
        30807 => X"63",  -- 99
        30808 => X"0C",  -- 12
        30809 => X"18",  -- 24
        30810 => X"63",  -- 99
        30811 => X"4F",  -- 79
        30812 => X"13",  -- 19
        30813 => X"5E",  -- 94
        30814 => X"55",  -- 85
        30815 => X"50",  -- 80
        30816 => X"64",  -- 100
        30817 => X"6E",  -- 110
        30818 => X"43",  -- 67
        30819 => X"0C",  -- 12
        30820 => X"23",  -- 35
        30821 => X"64",  -- 100
        30822 => X"42",  -- 66
        30823 => X"1F",  -- 31
        30824 => X"62",  -- 98
        30825 => X"22",  -- 34
        30826 => X"3E",  -- 62
        30827 => X"8E",  -- 142
        30828 => X"80",  -- 128
        30829 => X"3A",  -- 58
        30830 => X"99",  -- 153
        30831 => X"CE",  -- 206
        30832 => X"D9",  -- 217
        30833 => X"CF",  -- 207
        30834 => X"D4",  -- 212
        30835 => X"C3",  -- 195
        30836 => X"8A",  -- 138
        30837 => X"89",  -- 137
        30838 => X"92",  -- 146
        30839 => X"A0",  -- 160
        30840 => X"BD",  -- 189
        30841 => X"DD",  -- 221
        30842 => X"E3",  -- 227
        30843 => X"E3",  -- 227
        30844 => X"92",  -- 146
        30845 => X"22",  -- 34
        30846 => X"13",  -- 19
        30847 => X"1C",  -- 28
        30848 => X"5B",  -- 91
        30849 => X"8E",  -- 142
        30850 => X"99",  -- 153
        30851 => X"9A",  -- 154
        30852 => X"BD",  -- 189
        30853 => X"C3",  -- 195
        30854 => X"AF",  -- 175
        30855 => X"4B",  -- 75
        30856 => X"1E",  -- 30
        30857 => X"17",  -- 23
        30858 => X"0E",  -- 14
        30859 => X"1B",  -- 27
        30860 => X"51",  -- 81
        30861 => X"68",  -- 104
        30862 => X"96",  -- 150
        30863 => X"B7",  -- 183
        30864 => X"BF",  -- 191
        30865 => X"BC",  -- 188
        30866 => X"B6",  -- 182
        30867 => X"C4",  -- 196
        30868 => X"C0",  -- 192
        30869 => X"B4",  -- 180
        30870 => X"A4",  -- 164
        30871 => X"73",  -- 115
        30872 => X"36",  -- 54
        30873 => X"0B",  -- 11
        30874 => X"12",  -- 18
        30875 => X"12",  -- 18
        30876 => X"1E",  -- 30
        30877 => X"36",  -- 54
        30878 => X"72",  -- 114
        30879 => X"A1",  -- 161
        30880 => X"A7",  -- 167
        30881 => X"A7",  -- 167
        30882 => X"A7",  -- 167
        30883 => X"A5",  -- 165
        30884 => X"A7",  -- 167
        30885 => X"B0",  -- 176
        30886 => X"B9",  -- 185
        30887 => X"BE",  -- 190
        30888 => X"BE",  -- 190
        30889 => X"BC",  -- 188
        30890 => X"B9",  -- 185
        30891 => X"B8",  -- 184
        30892 => X"B8",  -- 184
        30893 => X"B2",  -- 178
        30894 => X"AA",  -- 170
        30895 => X"A5",  -- 165
        30896 => X"A6",  -- 166
        30897 => X"7B",  -- 123
        30898 => X"58",  -- 88
        30899 => X"4C",  -- 76
        30900 => X"36",  -- 54
        30901 => X"16",  -- 22
        30902 => X"0E",  -- 14
        30903 => X"1B",  -- 27
        30904 => X"24",  -- 36
        30905 => X"22",  -- 34
        30906 => X"17",  -- 23
        30907 => X"0E",  -- 14
        30908 => X"15",  -- 21
        30909 => X"32",  -- 50
        30910 => X"55",  -- 85
        30911 => X"6A",  -- 106
        30912 => X"7C",  -- 124
        30913 => X"6B",  -- 107
        30914 => X"68",  -- 104
        30915 => X"61",  -- 97
        30916 => X"49",  -- 73
        30917 => X"3E",  -- 62
        30918 => X"33",  -- 51
        30919 => X"19",  -- 25
        30920 => X"21",  -- 33
        30921 => X"2B",  -- 43
        30922 => X"43",  -- 67
        30923 => X"5E",  -- 94
        30924 => X"77",  -- 119
        30925 => X"8D",  -- 141
        30926 => X"A4",  -- 164
        30927 => X"B5",  -- 181
        30928 => X"BF",  -- 191
        30929 => X"B3",  -- 179
        30930 => X"B0",  -- 176
        30931 => X"B9",  -- 185
        30932 => X"C1",  -- 193
        30933 => X"BC",  -- 188
        30934 => X"B6",  -- 182
        30935 => X"B3",  -- 179
        30936 => X"BB",  -- 187
        30937 => X"B7",  -- 183
        30938 => X"B7",  -- 183
        30939 => X"BD",  -- 189
        30940 => X"C3",  -- 195
        30941 => X"BF",  -- 191
        30942 => X"B2",  -- 178
        30943 => X"A8",  -- 168
        30944 => X"9A",  -- 154
        30945 => X"7B",  -- 123
        30946 => X"76",  -- 118
        30947 => X"90",  -- 144
        30948 => X"A9",  -- 169
        30949 => X"B7",  -- 183
        30950 => X"C0",  -- 192
        30951 => X"C1",  -- 193
        30952 => X"C3",  -- 195
        30953 => X"C5",  -- 197
        30954 => X"C9",  -- 201
        30955 => X"CB",  -- 203
        30956 => X"C9",  -- 201
        30957 => X"C7",  -- 199
        30958 => X"C4",  -- 196
        30959 => X"C1",  -- 193
        30960 => X"B4",  -- 180
        30961 => X"AA",  -- 170
        30962 => X"AF",  -- 175
        30963 => X"9D",  -- 157
        30964 => X"78",  -- 120
        30965 => X"4F",  -- 79
        30966 => X"32",  -- 50
        30967 => X"37",  -- 55
        30968 => X"36",  -- 54
        30969 => X"29",  -- 41
        30970 => X"25",  -- 37
        30971 => X"40",  -- 64
        30972 => X"72",  -- 114
        30973 => X"95",  -- 149
        30974 => X"A9",  -- 169
        30975 => X"B8",  -- 184
        30976 => X"BE",  -- 190
        30977 => X"BA",  -- 186
        30978 => X"B8",  -- 184
        30979 => X"C3",  -- 195
        30980 => X"B1",  -- 177
        30981 => X"B2",  -- 178
        30982 => X"AA",  -- 170
        30983 => X"A8",  -- 168
        30984 => X"B4",  -- 180
        30985 => X"B9",  -- 185
        30986 => X"AE",  -- 174
        30987 => X"B5",  -- 181
        30988 => X"AC",  -- 172
        30989 => X"C4",  -- 196
        30990 => X"A2",  -- 162
        30991 => X"B6",  -- 182
        30992 => X"B0",  -- 176
        30993 => X"9E",  -- 158
        30994 => X"A8",  -- 168
        30995 => X"B0",  -- 176
        30996 => X"99",  -- 153
        30997 => X"B4",  -- 180
        30998 => X"B4",  -- 180
        30999 => X"A2",  -- 162
        31000 => X"9E",  -- 158
        31001 => X"9D",  -- 157
        31002 => X"9E",  -- 158
        31003 => X"8E",  -- 142
        31004 => X"8F",  -- 143
        31005 => X"8C",  -- 140
        31006 => X"7B",  -- 123
        31007 => X"8E",  -- 142
        31008 => X"98",  -- 152
        31009 => X"9A",  -- 154
        31010 => X"96",  -- 150
        31011 => X"91",  -- 145
        31012 => X"94",  -- 148
        31013 => X"9D",  -- 157
        31014 => X"9C",  -- 156
        31015 => X"95",  -- 149
        31016 => X"AD",  -- 173
        31017 => X"B5",  -- 181
        31018 => X"BA",  -- 186
        31019 => X"B7",  -- 183
        31020 => X"B5",  -- 181
        31021 => X"B7",  -- 183
        31022 => X"B6",  -- 182
        31023 => X"B0",  -- 176
        31024 => X"B1",  -- 177
        31025 => X"BD",  -- 189
        31026 => X"C4",  -- 196
        31027 => X"C0",  -- 192
        31028 => X"B8",  -- 184
        31029 => X"B7",  -- 183
        31030 => X"B8",  -- 184
        31031 => X"B8",  -- 184
        31032 => X"B6",  -- 182
        31033 => X"B6",  -- 182
        31034 => X"B7",  -- 183
        31035 => X"BC",  -- 188
        31036 => X"C3",  -- 195
        31037 => X"C4",  -- 196
        31038 => X"BC",  -- 188
        31039 => X"B0",  -- 176
        31040 => X"4F",  -- 79
        31041 => X"4E",  -- 78
        31042 => X"4D",  -- 77
        31043 => X"4F",  -- 79
        31044 => X"54",  -- 84
        31045 => X"5A",  -- 90
        31046 => X"5F",  -- 95
        31047 => X"63",  -- 99
        31048 => X"63",  -- 99
        31049 => X"60",  -- 96
        31050 => X"5C",  -- 92
        31051 => X"58",  -- 88
        31052 => X"54",  -- 84
        31053 => X"4F",  -- 79
        31054 => X"4C",  -- 76
        31055 => X"49",  -- 73
        31056 => X"49",  -- 73
        31057 => X"49",  -- 73
        31058 => X"4B",  -- 75
        31059 => X"4A",  -- 74
        31060 => X"48",  -- 72
        31061 => X"48",  -- 72
        31062 => X"46",  -- 70
        31063 => X"45",  -- 69
        31064 => X"44",  -- 68
        31065 => X"46",  -- 70
        31066 => X"49",  -- 73
        31067 => X"4E",  -- 78
        31068 => X"54",  -- 84
        31069 => X"57",  -- 87
        31070 => X"54",  -- 84
        31071 => X"4F",  -- 79
        31072 => X"5A",  -- 90
        31073 => X"75",  -- 117
        31074 => X"7B",  -- 123
        31075 => X"58",  -- 88
        31076 => X"2A",  -- 42
        31077 => X"10",  -- 16
        31078 => X"09",  -- 9
        31079 => X"08",  -- 8
        31080 => X"17",  -- 23
        31081 => X"3F",  -- 63
        31082 => X"6B",  -- 107
        31083 => X"7E",  -- 126
        31084 => X"82",  -- 130
        31085 => X"80",  -- 128
        31086 => X"7C",  -- 124
        31087 => X"84",  -- 132
        31088 => X"85",  -- 133
        31089 => X"84",  -- 132
        31090 => X"80",  -- 128
        31091 => X"6C",  -- 108
        31092 => X"42",  -- 66
        31093 => X"1D",  -- 29
        31094 => X"19",  -- 25
        31095 => X"29",  -- 41
        31096 => X"76",  -- 118
        31097 => X"95",  -- 149
        31098 => X"8A",  -- 138
        31099 => X"7E",  -- 126
        31100 => X"55",  -- 85
        31101 => X"2A",  -- 42
        31102 => X"35",  -- 53
        31103 => X"36",  -- 54
        31104 => X"1F",  -- 31
        31105 => X"5B",  -- 91
        31106 => X"BA",  -- 186
        31107 => X"BB",  -- 187
        31108 => X"A5",  -- 165
        31109 => X"8E",  -- 142
        31110 => X"94",  -- 148
        31111 => X"95",  -- 149
        31112 => X"B0",  -- 176
        31113 => X"CB",  -- 203
        31114 => X"E5",  -- 229
        31115 => X"D8",  -- 216
        31116 => X"D5",  -- 213
        31117 => X"DE",  -- 222
        31118 => X"96",  -- 150
        31119 => X"22",  -- 34
        31120 => X"48",  -- 72
        31121 => X"88",  -- 136
        31122 => X"6E",  -- 110
        31123 => X"41",  -- 65
        31124 => X"23",  -- 35
        31125 => X"4F",  -- 79
        31126 => X"6E",  -- 110
        31127 => X"42",  -- 66
        31128 => X"0F",  -- 15
        31129 => X"40",  -- 64
        31130 => X"77",  -- 119
        31131 => X"3A",  -- 58
        31132 => X"0C",  -- 12
        31133 => X"5E",  -- 94
        31134 => X"58",  -- 88
        31135 => X"41",  -- 65
        31136 => X"65",  -- 101
        31137 => X"77",  -- 119
        31138 => X"41",  -- 65
        31139 => X"1E",  -- 30
        31140 => X"1A",  -- 26
        31141 => X"6E",  -- 110
        31142 => X"46",  -- 70
        31143 => X"23",  -- 35
        31144 => X"64",  -- 100
        31145 => X"2A",  -- 42
        31146 => X"1A",  -- 26
        31147 => X"59",  -- 89
        31148 => X"69",  -- 105
        31149 => X"21",  -- 33
        31150 => X"7A",  -- 122
        31151 => X"C5",  -- 197
        31152 => X"CF",  -- 207
        31153 => X"D5",  -- 213
        31154 => X"D5",  -- 213
        31155 => X"B8",  -- 184
        31156 => X"83",  -- 131
        31157 => X"82",  -- 130
        31158 => X"7F",  -- 127
        31159 => X"8A",  -- 138
        31160 => X"BD",  -- 189
        31161 => X"DC",  -- 220
        31162 => X"DF",  -- 223
        31163 => X"E2",  -- 226
        31164 => X"B0",  -- 176
        31165 => X"43",  -- 67
        31166 => X"16",  -- 22
        31167 => X"1F",  -- 31
        31168 => X"26",  -- 38
        31169 => X"2E",  -- 46
        31170 => X"23",  -- 35
        31171 => X"28",  -- 40
        31172 => X"55",  -- 85
        31173 => X"81",  -- 129
        31174 => X"9D",  -- 157
        31175 => X"54",  -- 84
        31176 => X"17",  -- 23
        31177 => X"16",  -- 22
        31178 => X"1F",  -- 31
        31179 => X"3F",  -- 63
        31180 => X"85",  -- 133
        31181 => X"9E",  -- 158
        31182 => X"AE",  -- 174
        31183 => X"AF",  -- 175
        31184 => X"C1",  -- 193
        31185 => X"C2",  -- 194
        31186 => X"BD",  -- 189
        31187 => X"C9",  -- 201
        31188 => X"C2",  -- 194
        31189 => X"B9",  -- 185
        31190 => X"B5",  -- 181
        31191 => X"95",  -- 149
        31192 => X"50",  -- 80
        31193 => X"18",  -- 24
        31194 => X"14",  -- 20
        31195 => X"14",  -- 20
        31196 => X"24",  -- 36
        31197 => X"3E",  -- 62
        31198 => X"79",  -- 121
        31199 => X"AA",  -- 170
        31200 => X"B4",  -- 180
        31201 => X"B1",  -- 177
        31202 => X"A8",  -- 168
        31203 => X"A1",  -- 161
        31204 => X"A7",  -- 167
        31205 => X"B5",  -- 181
        31206 => X"BC",  -- 188
        31207 => X"B9",  -- 185
        31208 => X"C1",  -- 193
        31209 => X"BC",  -- 188
        31210 => X"B6",  -- 182
        31211 => X"B7",  -- 183
        31212 => X"BA",  -- 186
        31213 => X"BA",  -- 186
        31214 => X"B3",  -- 179
        31215 => X"AD",  -- 173
        31216 => X"9E",  -- 158
        31217 => X"9A",  -- 154
        31218 => X"85",  -- 133
        31219 => X"5F",  -- 95
        31220 => X"41",  -- 65
        31221 => X"32",  -- 50
        31222 => X"29",  -- 41
        31223 => X"20",  -- 32
        31224 => X"1F",  -- 31
        31225 => X"1B",  -- 27
        31226 => X"11",  -- 17
        31227 => X"0B",  -- 11
        31228 => X"1D",  -- 29
        31229 => X"41",  -- 65
        31230 => X"5F",  -- 95
        31231 => X"6C",  -- 108
        31232 => X"7A",  -- 122
        31233 => X"78",  -- 120
        31234 => X"6D",  -- 109
        31235 => X"5D",  -- 93
        31236 => X"4D",  -- 77
        31237 => X"3B",  -- 59
        31238 => X"30",  -- 48
        31239 => X"2E",  -- 46
        31240 => X"26",  -- 38
        31241 => X"31",  -- 49
        31242 => X"47",  -- 71
        31243 => X"62",  -- 98
        31244 => X"7B",  -- 123
        31245 => X"90",  -- 144
        31246 => X"A6",  -- 166
        31247 => X"B5",  -- 181
        31248 => X"C5",  -- 197
        31249 => X"BE",  -- 190
        31250 => X"BB",  -- 187
        31251 => X"BD",  -- 189
        31252 => X"C1",  -- 193
        31253 => X"C0",  -- 192
        31254 => X"BC",  -- 188
        31255 => X"BB",  -- 187
        31256 => X"AF",  -- 175
        31257 => X"AE",  -- 174
        31258 => X"B3",  -- 179
        31259 => X"BD",  -- 189
        31260 => X"C4",  -- 196
        31261 => X"C2",  -- 194
        31262 => X"B5",  -- 181
        31263 => X"AA",  -- 170
        31264 => X"97",  -- 151
        31265 => X"7D",  -- 125
        31266 => X"7D",  -- 125
        31267 => X"9B",  -- 155
        31268 => X"B2",  -- 178
        31269 => X"BC",  -- 188
        31270 => X"BE",  -- 190
        31271 => X"BA",  -- 186
        31272 => X"C2",  -- 194
        31273 => X"C8",  -- 200
        31274 => X"CC",  -- 204
        31275 => X"CE",  -- 206
        31276 => X"CD",  -- 205
        31277 => X"C7",  -- 199
        31278 => X"C1",  -- 193
        31279 => X"BD",  -- 189
        31280 => X"C0",  -- 192
        31281 => X"B3",  -- 179
        31282 => X"9F",  -- 159
        31283 => X"77",  -- 119
        31284 => X"5F",  -- 95
        31285 => X"58",  -- 88
        31286 => X"44",  -- 68
        31287 => X"3B",  -- 59
        31288 => X"36",  -- 54
        31289 => X"2F",  -- 47
        31290 => X"39",  -- 57
        31291 => X"57",  -- 87
        31292 => X"79",  -- 121
        31293 => X"94",  -- 148
        31294 => X"A3",  -- 163
        31295 => X"AD",  -- 173
        31296 => X"B1",  -- 177
        31297 => X"BF",  -- 191
        31298 => X"BB",  -- 187
        31299 => X"B1",  -- 177
        31300 => X"97",  -- 151
        31301 => X"A6",  -- 166
        31302 => X"AC",  -- 172
        31303 => X"AD",  -- 173
        31304 => X"9C",  -- 156
        31305 => X"B4",  -- 180
        31306 => X"B6",  -- 182
        31307 => X"AD",  -- 173
        31308 => X"A1",  -- 161
        31309 => X"B8",  -- 184
        31310 => X"A3",  -- 163
        31311 => X"B2",  -- 178
        31312 => X"AF",  -- 175
        31313 => X"9C",  -- 156
        31314 => X"A5",  -- 165
        31315 => X"AD",  -- 173
        31316 => X"96",  -- 150
        31317 => X"AD",  -- 173
        31318 => X"AC",  -- 172
        31319 => X"A0",  -- 160
        31320 => X"9F",  -- 159
        31321 => X"9A",  -- 154
        31322 => X"9C",  -- 156
        31323 => X"90",  -- 144
        31324 => X"90",  -- 144
        31325 => X"92",  -- 146
        31326 => X"7F",  -- 127
        31327 => X"81",  -- 129
        31328 => X"85",  -- 133
        31329 => X"87",  -- 135
        31330 => X"8E",  -- 142
        31331 => X"94",  -- 148
        31332 => X"9A",  -- 154
        31333 => X"9C",  -- 156
        31334 => X"A0",  -- 160
        31335 => X"A5",  -- 165
        31336 => X"AA",  -- 170
        31337 => X"B1",  -- 177
        31338 => X"B6",  -- 182
        31339 => X"B7",  -- 183
        31340 => X"B9",  -- 185
        31341 => X"BC",  -- 188
        31342 => X"B9",  -- 185
        31343 => X"B5",  -- 181
        31344 => X"B0",  -- 176
        31345 => X"BB",  -- 187
        31346 => X"C1",  -- 193
        31347 => X"BC",  -- 188
        31348 => X"B4",  -- 180
        31349 => X"B2",  -- 178
        31350 => X"B3",  -- 179
        31351 => X"B4",  -- 180
        31352 => X"B4",  -- 180
        31353 => X"B7",  -- 183
        31354 => X"BA",  -- 186
        31355 => X"BB",  -- 187
        31356 => X"BD",  -- 189
        31357 => X"BE",  -- 190
        31358 => X"B7",  -- 183
        31359 => X"AF",  -- 175
        31360 => X"50",  -- 80
        31361 => X"4F",  -- 79
        31362 => X"4D",  -- 77
        31363 => X"4D",  -- 77
        31364 => X"52",  -- 82
        31365 => X"58",  -- 88
        31366 => X"5E",  -- 94
        31367 => X"63",  -- 99
        31368 => X"66",  -- 102
        31369 => X"65",  -- 101
        31370 => X"64",  -- 100
        31371 => X"62",  -- 98
        31372 => X"5E",  -- 94
        31373 => X"57",  -- 87
        31374 => X"51",  -- 81
        31375 => X"4A",  -- 74
        31376 => X"4B",  -- 75
        31377 => X"4B",  -- 75
        31378 => X"4C",  -- 76
        31379 => X"4C",  -- 76
        31380 => X"4C",  -- 76
        31381 => X"4A",  -- 74
        31382 => X"49",  -- 73
        31383 => X"48",  -- 72
        31384 => X"47",  -- 71
        31385 => X"48",  -- 72
        31386 => X"4B",  -- 75
        31387 => X"4F",  -- 79
        31388 => X"51",  -- 81
        31389 => X"4E",  -- 78
        31390 => X"49",  -- 73
        31391 => X"45",  -- 69
        31392 => X"64",  -- 100
        31393 => X"81",  -- 129
        31394 => X"83",  -- 131
        31395 => X"56",  -- 86
        31396 => X"23",  -- 35
        31397 => X"0F",  -- 15
        31398 => X"0D",  -- 13
        31399 => X"0A",  -- 10
        31400 => X"1B",  -- 27
        31401 => X"49",  -- 73
        31402 => X"67",  -- 103
        31403 => X"71",  -- 113
        31404 => X"7F",  -- 127
        31405 => X"7C",  -- 124
        31406 => X"76",  -- 118
        31407 => X"83",  -- 131
        31408 => X"7A",  -- 122
        31409 => X"8A",  -- 138
        31410 => X"88",  -- 136
        31411 => X"62",  -- 98
        31412 => X"2E",  -- 46
        31413 => X"12",  -- 18
        31414 => X"19",  -- 25
        31415 => X"29",  -- 41
        31416 => X"68",  -- 104
        31417 => X"63",  -- 99
        31418 => X"3C",  -- 60
        31419 => X"31",  -- 49
        31420 => X"28",  -- 40
        31421 => X"16",  -- 22
        31422 => X"2C",  -- 44
        31423 => X"40",  -- 64
        31424 => X"29",  -- 41
        31425 => X"68",  -- 104
        31426 => X"BD",  -- 189
        31427 => X"B6",  -- 182
        31428 => X"A6",  -- 166
        31429 => X"7C",  -- 124
        31430 => X"91",  -- 145
        31431 => X"A8",  -- 168
        31432 => X"C2",  -- 194
        31433 => X"C8",  -- 200
        31434 => X"DA",  -- 218
        31435 => X"D3",  -- 211
        31436 => X"D8",  -- 216
        31437 => X"B7",  -- 183
        31438 => X"54",  -- 84
        31439 => X"21",  -- 33
        31440 => X"6B",  -- 107
        31441 => X"6F",  -- 111
        31442 => X"2A",  -- 42
        31443 => X"0D",  -- 13
        31444 => X"1A",  -- 26
        31445 => X"5F",  -- 95
        31446 => X"65",  -- 101
        31447 => X"23",  -- 35
        31448 => X"14",  -- 20
        31449 => X"5C",  -- 92
        31450 => X"75",  -- 117
        31451 => X"28",  -- 40
        31452 => X"0E",  -- 14
        31453 => X"4A",  -- 74
        31454 => X"4C",  -- 76
        31455 => X"3C",  -- 60
        31456 => X"60",  -- 96
        31457 => X"74",  -- 116
        31458 => X"4F",  -- 79
        31459 => X"28",  -- 40
        31460 => X"0C",  -- 12
        31461 => X"63",  -- 99
        31462 => X"57",  -- 87
        31463 => X"35",  -- 53
        31464 => X"75",  -- 117
        31465 => X"43",  -- 67
        31466 => X"09",  -- 9
        31467 => X"24",  -- 36
        31468 => X"5D",  -- 93
        31469 => X"17",  -- 23
        31470 => X"49",  -- 73
        31471 => X"AF",  -- 175
        31472 => X"BE",  -- 190
        31473 => X"CB",  -- 203
        31474 => X"D1",  -- 209
        31475 => X"C7",  -- 199
        31476 => X"A1",  -- 161
        31477 => X"92",  -- 146
        31478 => X"7D",  -- 125
        31479 => X"8F",  -- 143
        31480 => X"CE",  -- 206
        31481 => X"DC",  -- 220
        31482 => X"E1",  -- 225
        31483 => X"B9",  -- 185
        31484 => X"86",  -- 134
        31485 => X"7C",  -- 124
        31486 => X"61",  -- 97
        31487 => X"18",  -- 24
        31488 => X"14",  -- 20
        31489 => X"0C",  -- 12
        31490 => X"12",  -- 18
        31491 => X"1B",  -- 27
        31492 => X"29",  -- 41
        31493 => X"5F",  -- 95
        31494 => X"97",  -- 151
        31495 => X"68",  -- 104
        31496 => X"16",  -- 22
        31497 => X"0B",  -- 11
        31498 => X"14",  -- 20
        31499 => X"3A",  -- 58
        31500 => X"8E",  -- 142
        31501 => X"B5",  -- 181
        31502 => X"BE",  -- 190
        31503 => X"B4",  -- 180
        31504 => X"C3",  -- 195
        31505 => X"C4",  -- 196
        31506 => X"C0",  -- 192
        31507 => X"C6",  -- 198
        31508 => X"BF",  -- 191
        31509 => X"B4",  -- 180
        31510 => X"AF",  -- 175
        31511 => X"99",  -- 153
        31512 => X"67",  -- 103
        31513 => X"22",  -- 34
        31514 => X"12",  -- 18
        31515 => X"10",  -- 16
        31516 => X"1B",  -- 27
        31517 => X"2D",  -- 45
        31518 => X"68",  -- 104
        31519 => X"9D",  -- 157
        31520 => X"BB",  -- 187
        31521 => X"BA",  -- 186
        31522 => X"B0",  -- 176
        31523 => X"A4",  -- 164
        31524 => X"A6",  -- 166
        31525 => X"B6",  -- 182
        31526 => X"C0",  -- 192
        31527 => X"BF",  -- 191
        31528 => X"CD",  -- 205
        31529 => X"C4",  -- 196
        31530 => X"BB",  -- 187
        31531 => X"B8",  -- 184
        31532 => X"B9",  -- 185
        31533 => X"B9",  -- 185
        31534 => X"B2",  -- 178
        31535 => X"AA",  -- 170
        31536 => X"A5",  -- 165
        31537 => X"A4",  -- 164
        31538 => X"96",  -- 150
        31539 => X"7C",  -- 124
        31540 => X"5C",  -- 92
        31541 => X"40",  -- 64
        31542 => X"2F",  -- 47
        31543 => X"26",  -- 38
        31544 => X"21",  -- 33
        31545 => X"1F",  -- 31
        31546 => X"16",  -- 22
        31547 => X"15",  -- 21
        31548 => X"2F",  -- 47
        31549 => X"56",  -- 86
        31550 => X"6B",  -- 107
        31551 => X"6D",  -- 109
        31552 => X"69",  -- 105
        31553 => X"7A",  -- 122
        31554 => X"6F",  -- 111
        31555 => X"5C",  -- 92
        31556 => X"51",  -- 81
        31557 => X"35",  -- 53
        31558 => X"22",  -- 34
        31559 => X"2F",  -- 47
        31560 => X"30",  -- 48
        31561 => X"3B",  -- 59
        31562 => X"50",  -- 80
        31563 => X"68",  -- 104
        31564 => X"7D",  -- 125
        31565 => X"8F",  -- 143
        31566 => X"A1",  -- 161
        31567 => X"AD",  -- 173
        31568 => X"BE",  -- 190
        31569 => X"C1",  -- 193
        31570 => X"C2",  -- 194
        31571 => X"BE",  -- 190
        31572 => X"BC",  -- 188
        31573 => X"BC",  -- 188
        31574 => X"BA",  -- 186
        31575 => X"B9",  -- 185
        31576 => X"B6",  -- 182
        31577 => X"B0",  -- 176
        31578 => X"AC",  -- 172
        31579 => X"B0",  -- 176
        31580 => X"B9",  -- 185
        31581 => X"BE",  -- 190
        31582 => X"BB",  -- 187
        31583 => X"B5",  -- 181
        31584 => X"8E",  -- 142
        31585 => X"7B",  -- 123
        31586 => X"80",  -- 128
        31587 => X"A0",  -- 160
        31588 => X"B8",  -- 184
        31589 => X"C3",  -- 195
        31590 => X"C8",  -- 200
        31591 => X"C5",  -- 197
        31592 => X"C2",  -- 194
        31593 => X"C9",  -- 201
        31594 => X"CF",  -- 207
        31595 => X"D3",  -- 211
        31596 => X"CF",  -- 207
        31597 => X"C8",  -- 200
        31598 => X"C1",  -- 193
        31599 => X"BC",  -- 188
        31600 => X"AF",  -- 175
        31601 => X"B6",  -- 182
        31602 => X"AF",  -- 175
        31603 => X"7C",  -- 124
        31604 => X"52",  -- 82
        31605 => X"49",  -- 73
        31606 => X"43",  -- 67
        31607 => X"46",  -- 70
        31608 => X"32",  -- 50
        31609 => X"30",  -- 48
        31610 => X"4D",  -- 77
        31611 => X"70",  -- 112
        31612 => X"85",  -- 133
        31613 => X"9B",  -- 155
        31614 => X"B0",  -- 176
        31615 => X"B3",  -- 179
        31616 => X"A7",  -- 167
        31617 => X"BA",  -- 186
        31618 => X"B7",  -- 183
        31619 => X"B0",  -- 176
        31620 => X"9B",  -- 155
        31621 => X"A7",  -- 167
        31622 => X"A8",  -- 168
        31623 => X"AA",  -- 170
        31624 => X"97",  -- 151
        31625 => X"B5",  -- 181
        31626 => X"BF",  -- 191
        31627 => X"A7",  -- 167
        31628 => X"A1",  -- 161
        31629 => X"B2",  -- 178
        31630 => X"AB",  -- 171
        31631 => X"A9",  -- 169
        31632 => X"B0",  -- 176
        31633 => X"9B",  -- 155
        31634 => X"A4",  -- 164
        31635 => X"AD",  -- 173
        31636 => X"96",  -- 150
        31637 => X"A8",  -- 168
        31638 => X"A6",  -- 166
        31639 => X"A1",  -- 161
        31640 => X"98",  -- 152
        31641 => X"8E",  -- 142
        31642 => X"92",  -- 146
        31643 => X"8D",  -- 141
        31644 => X"8C",  -- 140
        31645 => X"94",  -- 148
        31646 => X"86",  -- 134
        31647 => X"77",  -- 119
        31648 => X"7C",  -- 124
        31649 => X"80",  -- 128
        31650 => X"8C",  -- 140
        31651 => X"98",  -- 152
        31652 => X"97",  -- 151
        31653 => X"93",  -- 147
        31654 => X"98",  -- 152
        31655 => X"A6",  -- 166
        31656 => X"B1",  -- 177
        31657 => X"B3",  -- 179
        31658 => X"B7",  -- 183
        31659 => X"B9",  -- 185
        31660 => X"BC",  -- 188
        31661 => X"BB",  -- 187
        31662 => X"B6",  -- 182
        31663 => X"AE",  -- 174
        31664 => X"AF",  -- 175
        31665 => X"B7",  -- 183
        31666 => X"BD",  -- 189
        31667 => X"BA",  -- 186
        31668 => X"B2",  -- 178
        31669 => X"B0",  -- 176
        31670 => X"B3",  -- 179
        31671 => X"B4",  -- 180
        31672 => X"B5",  -- 181
        31673 => X"BA",  -- 186
        31674 => X"BD",  -- 189
        31675 => X"BE",  -- 190
        31676 => X"BE",  -- 190
        31677 => X"BE",  -- 190
        31678 => X"B9",  -- 185
        31679 => X"B4",  -- 180
        31680 => X"53",  -- 83
        31681 => X"51",  -- 81
        31682 => X"4E",  -- 78
        31683 => X"4E",  -- 78
        31684 => X"52",  -- 82
        31685 => X"59",  -- 89
        31686 => X"5F",  -- 95
        31687 => X"64",  -- 100
        31688 => X"6A",  -- 106
        31689 => X"69",  -- 105
        31690 => X"68",  -- 104
        31691 => X"66",  -- 102
        31692 => X"63",  -- 99
        31693 => X"5C",  -- 92
        31694 => X"54",  -- 84
        31695 => X"4E",  -- 78
        31696 => X"4D",  -- 77
        31697 => X"4F",  -- 79
        31698 => X"53",  -- 83
        31699 => X"55",  -- 85
        31700 => X"55",  -- 85
        31701 => X"54",  -- 84
        31702 => X"52",  -- 82
        31703 => X"50",  -- 80
        31704 => X"4F",  -- 79
        31705 => X"4E",  -- 78
        31706 => X"51",  -- 81
        31707 => X"54",  -- 84
        31708 => X"54",  -- 84
        31709 => X"52",  -- 82
        31710 => X"4F",  -- 79
        31711 => X"50",  -- 80
        31712 => X"6E",  -- 110
        31713 => X"7F",  -- 127
        31714 => X"77",  -- 119
        31715 => X"4B",  -- 75
        31716 => X"1F",  -- 31
        31717 => X"0E",  -- 14
        31718 => X"0E",  -- 14
        31719 => X"0E",  -- 14
        31720 => X"22",  -- 34
        31721 => X"54",  -- 84
        31722 => X"54",  -- 84
        31723 => X"51",  -- 81
        31724 => X"6E",  -- 110
        31725 => X"77",  -- 119
        31726 => X"70",  -- 112
        31727 => X"74",  -- 116
        31728 => X"7E",  -- 126
        31729 => X"91",  -- 145
        31730 => X"92",  -- 146
        31731 => X"65",  -- 101
        31732 => X"2A",  -- 42
        31733 => X"13",  -- 19
        31734 => X"2B",  -- 43
        31735 => X"4E",  -- 78
        31736 => X"5A",  -- 90
        31737 => X"3D",  -- 61
        31738 => X"17",  -- 23
        31739 => X"14",  -- 20
        31740 => X"15",  -- 21
        31741 => X"14",  -- 20
        31742 => X"20",  -- 32
        31743 => X"12",  -- 18
        31744 => X"17",  -- 23
        31745 => X"51",  -- 81
        31746 => X"A0",  -- 160
        31747 => X"AA",  -- 170
        31748 => X"A4",  -- 164
        31749 => X"73",  -- 115
        31750 => X"6E",  -- 110
        31751 => X"AE",  -- 174
        31752 => X"C9",  -- 201
        31753 => X"DF",  -- 223
        31754 => X"D8",  -- 216
        31755 => X"D1",  -- 209
        31756 => X"D2",  -- 210
        31757 => X"80",  -- 128
        31758 => X"2F",  -- 47
        31759 => X"51",  -- 81
        31760 => X"6B",  -- 107
        31761 => X"2F",  -- 47
        31762 => X"0A",  -- 10
        31763 => X"11",  -- 17
        31764 => X"59",  -- 89
        31765 => X"72",  -- 114
        31766 => X"58",  -- 88
        31767 => X"0B",  -- 11
        31768 => X"1D",  -- 29
        31769 => X"5E",  -- 94
        31770 => X"5D",  -- 93
        31771 => X"18",  -- 24
        31772 => X"1B",  -- 27
        31773 => X"47",  -- 71
        31774 => X"4D",  -- 77
        31775 => X"3D",  -- 61
        31776 => X"58",  -- 88
        31777 => X"6E",  -- 110
        31778 => X"68",  -- 104
        31779 => X"2D",  -- 45
        31780 => X"09",  -- 9
        31781 => X"49",  -- 73
        31782 => X"6E",  -- 110
        31783 => X"50",  -- 80
        31784 => X"8B",  -- 139
        31785 => X"6D",  -- 109
        31786 => X"1A",  -- 26
        31787 => X"0E",  -- 14
        31788 => X"61",  -- 97
        31789 => X"36",  -- 54
        31790 => X"2A",  -- 42
        31791 => X"88",  -- 136
        31792 => X"C3",  -- 195
        31793 => X"C3",  -- 195
        31794 => X"C2",  -- 194
        31795 => X"C9",  -- 201
        31796 => X"B0",  -- 176
        31797 => X"87",  -- 135
        31798 => X"61",  -- 97
        31799 => X"82",  -- 130
        31800 => X"BA",  -- 186
        31801 => X"CF",  -- 207
        31802 => X"C8",  -- 200
        31803 => X"7F",  -- 127
        31804 => X"72",  -- 114
        31805 => X"C0",  -- 192
        31806 => X"AE",  -- 174
        31807 => X"39",  -- 57
        31808 => X"19",  -- 25
        31809 => X"0C",  -- 12
        31810 => X"1C",  -- 28
        31811 => X"1F",  -- 31
        31812 => X"13",  -- 19
        31813 => X"52",  -- 82
        31814 => X"9E",  -- 158
        31815 => X"7D",  -- 125
        31816 => X"31",  -- 49
        31817 => X"10",  -- 16
        31818 => X"14",  -- 20
        31819 => X"3A",  -- 58
        31820 => X"8B",  -- 139
        31821 => X"B4",  -- 180
        31822 => X"C3",  -- 195
        31823 => X"C2",  -- 194
        31824 => X"C6",  -- 198
        31825 => X"C5",  -- 197
        31826 => X"C4",  -- 196
        31827 => X"C8",  -- 200
        31828 => X"C3",  -- 195
        31829 => X"B7",  -- 183
        31830 => X"AA",  -- 170
        31831 => X"9C",  -- 156
        31832 => X"66",  -- 102
        31833 => X"22",  -- 34
        31834 => X"17",  -- 23
        31835 => X"1B",  -- 27
        31836 => X"25",  -- 37
        31837 => X"34",  -- 52
        31838 => X"70",  -- 112
        31839 => X"AD",  -- 173
        31840 => X"B4",  -- 180
        31841 => X"B6",  -- 182
        31842 => X"B3",  -- 179
        31843 => X"AC",  -- 172
        31844 => X"A7",  -- 167
        31845 => X"AC",  -- 172
        31846 => X"B9",  -- 185
        31847 => X"C4",  -- 196
        31848 => X"CE",  -- 206
        31849 => X"C7",  -- 199
        31850 => X"BF",  -- 191
        31851 => X"BA",  -- 186
        31852 => X"B7",  -- 183
        31853 => X"B3",  -- 179
        31854 => X"AD",  -- 173
        31855 => X"A8",  -- 168
        31856 => X"AB",  -- 171
        31857 => X"9D",  -- 157
        31858 => X"90",  -- 144
        31859 => X"87",  -- 135
        31860 => X"71",  -- 113
        31861 => X"4E",  -- 78
        31862 => X"32",  -- 50
        31863 => X"27",  -- 39
        31864 => X"21",  -- 33
        31865 => X"20",  -- 32
        31866 => X"1A",  -- 26
        31867 => X"1E",  -- 30
        31868 => X"3D",  -- 61
        31869 => X"66",  -- 102
        31870 => X"79",  -- 121
        31871 => X"77",  -- 119
        31872 => X"60",  -- 96
        31873 => X"6D",  -- 109
        31874 => X"6D",  -- 109
        31875 => X"66",  -- 102
        31876 => X"58",  -- 88
        31877 => X"39",  -- 57
        31878 => X"20",  -- 32
        31879 => X"20",  -- 32
        31880 => X"2D",  -- 45
        31881 => X"3A",  -- 58
        31882 => X"50",  -- 80
        31883 => X"68",  -- 104
        31884 => X"7C",  -- 124
        31885 => X"8E",  -- 142
        31886 => X"9E",  -- 158
        31887 => X"A8",  -- 168
        31888 => X"B0",  -- 176
        31889 => X"BC",  -- 188
        31890 => X"C4",  -- 196
        31891 => X"BF",  -- 191
        31892 => X"B8",  -- 184
        31893 => X"B7",  -- 183
        31894 => X"B6",  -- 182
        31895 => X"B3",  -- 179
        31896 => X"B9",  -- 185
        31897 => X"B2",  -- 178
        31898 => X"AB",  -- 171
        31899 => X"A9",  -- 169
        31900 => X"B0",  -- 176
        31901 => X"B7",  -- 183
        31902 => X"B5",  -- 181
        31903 => X"AE",  -- 174
        31904 => X"A1",  -- 161
        31905 => X"8D",  -- 141
        31906 => X"90",  -- 144
        31907 => X"A4",  -- 164
        31908 => X"B3",  -- 179
        31909 => X"B8",  -- 184
        31910 => X"BD",  -- 189
        31911 => X"BC",  -- 188
        31912 => X"C1",  -- 193
        31913 => X"C5",  -- 197
        31914 => X"CD",  -- 205
        31915 => X"D1",  -- 209
        31916 => X"CF",  -- 207
        31917 => X"C9",  -- 201
        31918 => X"C4",  -- 196
        31919 => X"C0",  -- 192
        31920 => X"BB",  -- 187
        31921 => X"AB",  -- 171
        31922 => X"9C",  -- 156
        31923 => X"7B",  -- 123
        31924 => X"60",  -- 96
        31925 => X"4E",  -- 78
        31926 => X"37",  -- 55
        31927 => X"30",  -- 48
        31928 => X"30",  -- 48
        31929 => X"2F",  -- 47
        31930 => X"55",  -- 85
        31931 => X"7D",  -- 125
        31932 => X"8B",  -- 139
        31933 => X"A1",  -- 161
        31934 => X"BA",  -- 186
        31935 => X"BB",  -- 187
        31936 => X"AC",  -- 172
        31937 => X"A9",  -- 169
        31938 => X"9F",  -- 159
        31939 => X"AE",  -- 174
        31940 => X"AF",  -- 175
        31941 => X"B0",  -- 176
        31942 => X"A5",  -- 165
        31943 => X"AD",  -- 173
        31944 => X"A5",  -- 165
        31945 => X"B3",  -- 179
        31946 => X"BC",  -- 188
        31947 => X"A2",  -- 162
        31948 => X"A8",  -- 168
        31949 => X"AF",  -- 175
        31950 => X"B0",  -- 176
        31951 => X"A2",  -- 162
        31952 => X"B0",  -- 176
        31953 => X"A0",  -- 160
        31954 => X"A7",  -- 167
        31955 => X"B0",  -- 176
        31956 => X"9C",  -- 156
        31957 => X"A7",  -- 167
        31958 => X"A0",  -- 160
        31959 => X"A0",  -- 160
        31960 => X"8D",  -- 141
        31961 => X"86",  -- 134
        31962 => X"8A",  -- 138
        31963 => X"86",  -- 134
        31964 => X"81",  -- 129
        31965 => X"8B",  -- 139
        31966 => X"8B",  -- 139
        31967 => X"79",  -- 121
        31968 => X"7D",  -- 125
        31969 => X"84",  -- 132
        31970 => X"8D",  -- 141
        31971 => X"94",  -- 148
        31972 => X"91",  -- 145
        31973 => X"8C",  -- 140
        31974 => X"93",  -- 147
        31975 => X"9E",  -- 158
        31976 => X"B1",  -- 177
        31977 => X"B1",  -- 177
        31978 => X"B4",  -- 180
        31979 => X"BA",  -- 186
        31980 => X"BC",  -- 188
        31981 => X"B9",  -- 185
        31982 => X"B0",  -- 176
        31983 => X"AB",  -- 171
        31984 => X"B1",  -- 177
        31985 => X"B8",  -- 184
        31986 => X"BE",  -- 190
        31987 => X"BB",  -- 187
        31988 => X"B7",  -- 183
        31989 => X"B6",  -- 182
        31990 => X"B7",  -- 183
        31991 => X"B7",  -- 183
        31992 => X"B5",  -- 181
        31993 => X"BA",  -- 186
        31994 => X"BE",  -- 190
        31995 => X"BE",  -- 190
        31996 => X"C1",  -- 193
        31997 => X"C0",  -- 192
        31998 => X"BB",  -- 187
        31999 => X"B4",  -- 180
        32000 => X"53",  -- 83
        32001 => X"51",  -- 81
        32002 => X"4E",  -- 78
        32003 => X"4E",  -- 78
        32004 => X"53",  -- 83
        32005 => X"59",  -- 89
        32006 => X"5F",  -- 95
        32007 => X"64",  -- 100
        32008 => X"67",  -- 103
        32009 => X"64",  -- 100
        32010 => X"60",  -- 96
        32011 => X"5E",  -- 94
        32012 => X"5B",  -- 91
        32013 => X"57",  -- 87
        32014 => X"50",  -- 80
        32015 => X"4B",  -- 75
        32016 => X"4C",  -- 76
        32017 => X"4F",  -- 79
        32018 => X"53",  -- 83
        32019 => X"58",  -- 88
        32020 => X"5A",  -- 90
        32021 => X"58",  -- 88
        32022 => X"56",  -- 86
        32023 => X"53",  -- 83
        32024 => X"56",  -- 86
        32025 => X"54",  -- 84
        32026 => X"56",  -- 86
        32027 => X"58",  -- 88
        32028 => X"55",  -- 85
        32029 => X"54",  -- 84
        32030 => X"56",  -- 86
        32031 => X"5E",  -- 94
        32032 => X"74",  -- 116
        32033 => X"71",  -- 113
        32034 => X"5F",  -- 95
        32035 => X"3D",  -- 61
        32036 => X"1B",  -- 27
        32037 => X"0C",  -- 12
        32038 => X"0A",  -- 10
        32039 => X"0B",  -- 11
        32040 => X"27",  -- 39
        32041 => X"62",  -- 98
        32042 => X"49",  -- 73
        32043 => X"2B",  -- 43
        32044 => X"45",  -- 69
        32045 => X"55",  -- 85
        32046 => X"56",  -- 86
        32047 => X"56",  -- 86
        32048 => X"64",  -- 100
        32049 => X"7A",  -- 122
        32050 => X"82",  -- 130
        32051 => X"59",  -- 89
        32052 => X"1A",  -- 26
        32053 => X"06",  -- 6
        32054 => X"3B",  -- 59
        32055 => X"7E",  -- 126
        32056 => X"6C",  -- 108
        32057 => X"33",  -- 51
        32058 => X"19",  -- 25
        32059 => X"20",  -- 32
        32060 => X"19",  -- 25
        32061 => X"2A",  -- 42
        32062 => X"4A",  -- 74
        32063 => X"3D",  -- 61
        32064 => X"1B",  -- 27
        32065 => X"30",  -- 48
        32066 => X"7D",  -- 125
        32067 => X"99",  -- 153
        32068 => X"7B",  -- 123
        32069 => X"75",  -- 117
        32070 => X"65",  -- 101
        32071 => X"A4",  -- 164
        32072 => X"A3",  -- 163
        32073 => X"DA",  -- 218
        32074 => X"D8",  -- 216
        32075 => X"D2",  -- 210
        32076 => X"C5",  -- 197
        32077 => X"85",  -- 133
        32078 => X"59",  -- 89
        32079 => X"5C",  -- 92
        32080 => X"44",  -- 68
        32081 => X"10",  -- 16
        32082 => X"0D",  -- 13
        32083 => X"3F",  -- 63
        32084 => X"83",  -- 131
        32085 => X"6E",  -- 110
        32086 => X"43",  -- 67
        32087 => X"0C",  -- 12
        32088 => X"38",  -- 56
        32089 => X"50",  -- 80
        32090 => X"3A",  -- 58
        32091 => X"1B",  -- 27
        32092 => X"39",  -- 57
        32093 => X"5F",  -- 95
        32094 => X"5A",  -- 90
        32095 => X"3E",  -- 62
        32096 => X"58",  -- 88
        32097 => X"6C",  -- 108
        32098 => X"6D",  -- 109
        32099 => X"3D",  -- 61
        32100 => X"0B",  -- 11
        32101 => X"43",  -- 67
        32102 => X"73",  -- 115
        32103 => X"50",  -- 80
        32104 => X"82",  -- 130
        32105 => X"8E",  -- 142
        32106 => X"55",  -- 85
        32107 => X"0C",  -- 12
        32108 => X"53",  -- 83
        32109 => X"69",  -- 105
        32110 => X"2E",  -- 46
        32111 => X"5E",  -- 94
        32112 => X"C3",  -- 195
        32113 => X"BF",  -- 191
        32114 => X"B4",  -- 180
        32115 => X"BC",  -- 188
        32116 => X"B1",  -- 177
        32117 => X"90",  -- 144
        32118 => X"68",  -- 104
        32119 => X"86",  -- 134
        32120 => X"B2",  -- 178
        32121 => X"D8",  -- 216
        32122 => X"BB",  -- 187
        32123 => X"89",  -- 137
        32124 => X"B5",  -- 181
        32125 => X"DB",  -- 219
        32126 => X"96",  -- 150
        32127 => X"4F",  -- 79
        32128 => X"24",  -- 36
        32129 => X"0D",  -- 13
        32130 => X"11",  -- 17
        32131 => X"14",  -- 20
        32132 => X"12",  -- 18
        32133 => X"73",  -- 115
        32134 => X"CA",  -- 202
        32135 => X"B1",  -- 177
        32136 => X"45",  -- 69
        32137 => X"13",  -- 19
        32138 => X"1F",  -- 31
        32139 => X"53",  -- 83
        32140 => X"A1",  -- 161
        32141 => X"BD",  -- 189
        32142 => X"BB",  -- 187
        32143 => X"BB",  -- 187
        32144 => X"B7",  -- 183
        32145 => X"B9",  -- 185
        32146 => X"B9",  -- 185
        32147 => X"B3",  -- 179
        32148 => X"A5",  -- 165
        32149 => X"97",  -- 151
        32150 => X"91",  -- 145
        32151 => X"9B",  -- 155
        32152 => X"54",  -- 84
        32153 => X"15",  -- 21
        32154 => X"11",  -- 17
        32155 => X"16",  -- 22
        32156 => X"1A",  -- 26
        32157 => X"22",  -- 34
        32158 => X"5C",  -- 92
        32159 => X"9B",  -- 155
        32160 => X"B2",  -- 178
        32161 => X"AD",  -- 173
        32162 => X"AC",  -- 172
        32163 => X"B2",  -- 178
        32164 => X"B0",  -- 176
        32165 => X"AB",  -- 171
        32166 => X"B0",  -- 176
        32167 => X"BB",  -- 187
        32168 => X"C1",  -- 193
        32169 => X"C2",  -- 194
        32170 => X"C1",  -- 193
        32171 => X"BC",  -- 188
        32172 => X"B5",  -- 181
        32173 => X"AF",  -- 175
        32174 => X"AA",  -- 170
        32175 => X"A9",  -- 169
        32176 => X"9E",  -- 158
        32177 => X"A0",  -- 160
        32178 => X"98",  -- 152
        32179 => X"88",  -- 136
        32180 => X"78",  -- 120
        32181 => X"67",  -- 103
        32182 => X"4D",  -- 77
        32183 => X"33",  -- 51
        32184 => X"23",  -- 35
        32185 => X"1E",  -- 30
        32186 => X"16",  -- 22
        32187 => X"1B",  -- 27
        32188 => X"3A",  -- 58
        32189 => X"65",  -- 101
        32190 => X"80",  -- 128
        32191 => X"86",  -- 134
        32192 => X"71",  -- 113
        32193 => X"64",  -- 100
        32194 => X"68",  -- 104
        32195 => X"6B",  -- 107
        32196 => X"5A",  -- 90
        32197 => X"48",  -- 72
        32198 => X"39",  -- 57
        32199 => X"26",  -- 38
        32200 => X"20",  -- 32
        32201 => X"31",  -- 49
        32202 => X"4B",  -- 75
        32203 => X"65",  -- 101
        32204 => X"7B",  -- 123
        32205 => X"90",  -- 144
        32206 => X"A0",  -- 160
        32207 => X"A8",  -- 168
        32208 => X"AC",  -- 172
        32209 => X"BA",  -- 186
        32210 => X"C2",  -- 194
        32211 => X"BB",  -- 187
        32212 => X"B4",  -- 180
        32213 => X"B5",  -- 181
        32214 => X"B7",  -- 183
        32215 => X"B8",  -- 184
        32216 => X"AE",  -- 174
        32217 => X"AF",  -- 175
        32218 => X"B1",  -- 177
        32219 => X"B4",  -- 180
        32220 => X"B8",  -- 184
        32221 => X"B7",  -- 183
        32222 => X"A9",  -- 169
        32223 => X"98",  -- 152
        32224 => X"98",  -- 152
        32225 => X"8B",  -- 139
        32226 => X"91",  -- 145
        32227 => X"A5",  -- 165
        32228 => X"B0",  -- 176
        32229 => X"B6",  -- 182
        32230 => X"BB",  -- 187
        32231 => X"BB",  -- 187
        32232 => X"BB",  -- 187
        32233 => X"BF",  -- 191
        32234 => X"C5",  -- 197
        32235 => X"C7",  -- 199
        32236 => X"C7",  -- 199
        32237 => X"C6",  -- 198
        32238 => X"C4",  -- 196
        32239 => X"C3",  -- 195
        32240 => X"C4",  -- 196
        32241 => X"AD",  -- 173
        32242 => X"95",  -- 149
        32243 => X"72",  -- 114
        32244 => X"5B",  -- 91
        32245 => X"4E",  -- 78
        32246 => X"37",  -- 55
        32247 => X"31",  -- 49
        32248 => X"36",  -- 54
        32249 => X"37",  -- 55
        32250 => X"5E",  -- 94
        32251 => X"86",  -- 134
        32252 => X"8F",  -- 143
        32253 => X"9E",  -- 158
        32254 => X"AF",  -- 175
        32255 => X"AA",  -- 170
        32256 => X"AC",  -- 172
        32257 => X"A2",  -- 162
        32258 => X"8E",  -- 142
        32259 => X"9E",  -- 158
        32260 => X"A9",  -- 169
        32261 => X"B3",  -- 179
        32262 => X"AB",  -- 171
        32263 => X"B9",  -- 185
        32264 => X"AE",  -- 174
        32265 => X"AE",  -- 174
        32266 => X"B4",  -- 180
        32267 => X"A4",  -- 164
        32268 => X"AB",  -- 171
        32269 => X"A3",  -- 163
        32270 => X"B2",  -- 178
        32271 => X"A8",  -- 168
        32272 => X"B5",  -- 181
        32273 => X"A7",  -- 167
        32274 => X"AB",  -- 171
        32275 => X"B0",  -- 176
        32276 => X"9D",  -- 157
        32277 => X"A5",  -- 165
        32278 => X"98",  -- 152
        32279 => X"96",  -- 150
        32280 => X"87",  -- 135
        32281 => X"84",  -- 132
        32282 => X"86",  -- 134
        32283 => X"82",  -- 130
        32284 => X"75",  -- 117
        32285 => X"7B",  -- 123
        32286 => X"8B",  -- 139
        32287 => X"84",  -- 132
        32288 => X"82",  -- 130
        32289 => X"8B",  -- 139
        32290 => X"90",  -- 144
        32291 => X"8E",  -- 142
        32292 => X"8E",  -- 142
        32293 => X"95",  -- 149
        32294 => X"9D",  -- 157
        32295 => X"A0",  -- 160
        32296 => X"AE",  -- 174
        32297 => X"AD",  -- 173
        32298 => X"B2",  -- 178
        32299 => X"BB",  -- 187
        32300 => X"BD",  -- 189
        32301 => X"B7",  -- 183
        32302 => X"B3",  -- 179
        32303 => X"B3",  -- 179
        32304 => X"B6",  -- 182
        32305 => X"BE",  -- 190
        32306 => X"C3",  -- 195
        32307 => X"C0",  -- 192
        32308 => X"BA",  -- 186
        32309 => X"B8",  -- 184
        32310 => X"B9",  -- 185
        32311 => X"B8",  -- 184
        32312 => X"B8",  -- 184
        32313 => X"B8",  -- 184
        32314 => X"B9",  -- 185
        32315 => X"BA",  -- 186
        32316 => X"BE",  -- 190
        32317 => X"BF",  -- 191
        32318 => X"B4",  -- 180
        32319 => X"A8",  -- 168
        32320 => X"57",  -- 87
        32321 => X"56",  -- 86
        32322 => X"54",  -- 84
        32323 => X"55",  -- 85
        32324 => X"59",  -- 89
        32325 => X"60",  -- 96
        32326 => X"65",  -- 101
        32327 => X"6A",  -- 106
        32328 => X"67",  -- 103
        32329 => X"62",  -- 98
        32330 => X"5C",  -- 92
        32331 => X"59",  -- 89
        32332 => X"58",  -- 88
        32333 => X"55",  -- 85
        32334 => X"51",  -- 81
        32335 => X"4C",  -- 76
        32336 => X"4C",  -- 76
        32337 => X"4F",  -- 79
        32338 => X"54",  -- 84
        32339 => X"58",  -- 88
        32340 => X"59",  -- 89
        32341 => X"58",  -- 88
        32342 => X"57",  -- 87
        32343 => X"55",  -- 85
        32344 => X"58",  -- 88
        32345 => X"56",  -- 86
        32346 => X"54",  -- 84
        32347 => X"55",  -- 85
        32348 => X"53",  -- 83
        32349 => X"52",  -- 82
        32350 => X"5A",  -- 90
        32351 => X"65",  -- 101
        32352 => X"7B",  -- 123
        32353 => X"6C",  -- 108
        32354 => X"53",  -- 83
        32355 => X"34",  -- 52
        32356 => X"1A",  -- 26
        32357 => X"0C",  -- 12
        32358 => X"09",  -- 9
        32359 => X"0A",  -- 10
        32360 => X"34",  -- 52
        32361 => X"72",  -- 114
        32362 => X"4E",  -- 78
        32363 => X"1B",  -- 27
        32364 => X"1E",  -- 30
        32365 => X"29",  -- 41
        32366 => X"37",  -- 55
        32367 => X"39",  -- 57
        32368 => X"57",  -- 87
        32369 => X"6C",  -- 108
        32370 => X"78",  -- 120
        32371 => X"57",  -- 87
        32372 => X"1C",  -- 28
        32373 => X"10",  -- 16
        32374 => X"59",  -- 89
        32375 => X"B4",  -- 180
        32376 => X"8A",  -- 138
        32377 => X"38",  -- 56
        32378 => X"19",  -- 25
        32379 => X"20",  -- 32
        32380 => X"19",  -- 25
        32381 => X"3E",  -- 62
        32382 => X"8D",  -- 141
        32383 => X"BA",  -- 186
        32384 => X"64",  -- 100
        32385 => X"1B",  -- 27
        32386 => X"45",  -- 69
        32387 => X"8B",  -- 139
        32388 => X"64",  -- 100
        32389 => X"7D",  -- 125
        32390 => X"83",  -- 131
        32391 => X"A3",  -- 163
        32392 => X"AA",  -- 170
        32393 => X"C1",  -- 193
        32394 => X"C9",  -- 201
        32395 => X"D2",  -- 210
        32396 => X"B3",  -- 179
        32397 => X"8E",  -- 142
        32398 => X"7A",  -- 122
        32399 => X"46",  -- 70
        32400 => X"2E",  -- 46
        32401 => X"28",  -- 40
        32402 => X"3A",  -- 58
        32403 => X"75",  -- 117
        32404 => X"7B",  -- 123
        32405 => X"70",  -- 112
        32406 => X"49",  -- 73
        32407 => X"38",  -- 56
        32408 => X"5C",  -- 92
        32409 => X"28",  -- 40
        32410 => X"1A",  -- 26
        32411 => X"40",  -- 64
        32412 => X"56",  -- 86
        32413 => X"60",  -- 96
        32414 => X"55",  -- 85
        32415 => X"4A",  -- 74
        32416 => X"59",  -- 89
        32417 => X"67",  -- 103
        32418 => X"53",  -- 83
        32419 => X"4A",  -- 74
        32420 => X"0B",  -- 11
        32421 => X"4D",  -- 77
        32422 => X"5D",  -- 93
        32423 => X"31",  -- 49
        32424 => X"58",  -- 88
        32425 => X"8A",  -- 138
        32426 => X"83",  -- 131
        32427 => X"18",  -- 24
        32428 => X"34",  -- 52
        32429 => X"79",  -- 121
        32430 => X"48",  -- 72
        32431 => X"46",  -- 70
        32432 => X"A5",  -- 165
        32433 => X"BA",  -- 186
        32434 => X"BE",  -- 190
        32435 => X"C2",  -- 194
        32436 => X"C3",  -- 195
        32437 => X"BA",  -- 186
        32438 => X"8C",  -- 140
        32439 => X"8C",  -- 140
        32440 => X"C3",  -- 195
        32441 => X"E0",  -- 224
        32442 => X"CF",  -- 207
        32443 => X"C3",  -- 195
        32444 => X"E3",  -- 227
        32445 => X"D9",  -- 217
        32446 => X"92",  -- 146
        32447 => X"54",  -- 84
        32448 => X"15",  -- 21
        32449 => X"22",  -- 34
        32450 => X"44",  -- 68
        32451 => X"56",  -- 86
        32452 => X"55",  -- 85
        32453 => X"A0",  -- 160
        32454 => X"CF",  -- 207
        32455 => X"B7",  -- 183
        32456 => X"56",  -- 86
        32457 => X"15",  -- 21
        32458 => X"27",  -- 39
        32459 => X"5E",  -- 94
        32460 => X"A8",  -- 168
        32461 => X"BE",  -- 190
        32462 => X"B6",  -- 182
        32463 => X"B8",  -- 184
        32464 => X"B8",  -- 184
        32465 => X"B6",  -- 182
        32466 => X"AC",  -- 172
        32467 => X"88",  -- 136
        32468 => X"63",  -- 99
        32469 => X"51",  -- 81
        32470 => X"5F",  -- 95
        32471 => X"8A",  -- 138
        32472 => X"64",  -- 100
        32473 => X"24",  -- 36
        32474 => X"1D",  -- 29
        32475 => X"20",  -- 32
        32476 => X"23",  -- 35
        32477 => X"2A",  -- 42
        32478 => X"60",  -- 96
        32479 => X"9A",  -- 154
        32480 => X"C1",  -- 193
        32481 => X"B1",  -- 177
        32482 => X"AB",  -- 171
        32483 => X"B3",  -- 179
        32484 => X"BA",  -- 186
        32485 => X"B6",  -- 182
        32486 => X"B3",  -- 179
        32487 => X"B3",  -- 179
        32488 => X"BD",  -- 189
        32489 => X"C2",  -- 194
        32490 => X"C4",  -- 196
        32491 => X"BE",  -- 190
        32492 => X"B2",  -- 178
        32493 => X"A8",  -- 168
        32494 => X"A2",  -- 162
        32495 => X"A2",  -- 162
        32496 => X"9A",  -- 154
        32497 => X"9A",  -- 154
        32498 => X"98",  -- 152
        32499 => X"91",  -- 145
        32500 => X"82",  -- 130
        32501 => X"6E",  -- 110
        32502 => X"5D",  -- 93
        32503 => X"53",  -- 83
        32504 => X"3C",  -- 60
        32505 => X"2B",  -- 43
        32506 => X"1B",  -- 27
        32507 => X"1D",  -- 29
        32508 => X"37",  -- 55
        32509 => X"5C",  -- 92
        32510 => X"7A",  -- 122
        32511 => X"89",  -- 137
        32512 => X"84",  -- 132
        32513 => X"63",  -- 99
        32514 => X"5C",  -- 92
        32515 => X"5F",  -- 95
        32516 => X"50",  -- 80
        32517 => X"4C",  -- 76
        32518 => X"4C",  -- 76
        32519 => X"39",  -- 57
        32520 => X"21",  -- 33
        32521 => X"35",  -- 53
        32522 => X"4F",  -- 79
        32523 => X"67",  -- 103
        32524 => X"7E",  -- 126
        32525 => X"90",  -- 144
        32526 => X"9E",  -- 158
        32527 => X"A3",  -- 163
        32528 => X"AE",  -- 174
        32529 => X"B4",  -- 180
        32530 => X"B7",  -- 183
        32531 => X"B1",  -- 177
        32532 => X"AC",  -- 172
        32533 => X"AF",  -- 175
        32534 => X"B6",  -- 182
        32535 => X"BD",  -- 189
        32536 => X"B4",  -- 180
        32537 => X"B6",  -- 182
        32538 => X"B7",  -- 183
        32539 => X"B7",  -- 183
        32540 => X"BC",  -- 188
        32541 => X"BC",  -- 188
        32542 => X"AF",  -- 175
        32543 => X"9E",  -- 158
        32544 => X"7D",  -- 125
        32545 => X"7A",  -- 122
        32546 => X"8A",  -- 138
        32547 => X"A4",  -- 164
        32548 => X"B3",  -- 179
        32549 => X"BC",  -- 188
        32550 => X"C6",  -- 198
        32551 => X"C8",  -- 200
        32552 => X"B7",  -- 183
        32553 => X"BA",  -- 186
        32554 => X"BC",  -- 188
        32555 => X"BE",  -- 190
        32556 => X"BF",  -- 191
        32557 => X"BF",  -- 191
        32558 => X"C0",  -- 192
        32559 => X"C2",  -- 194
        32560 => X"B6",  -- 182
        32561 => X"B4",  -- 180
        32562 => X"A4",  -- 164
        32563 => X"73",  -- 115
        32564 => X"53",  -- 83
        32565 => X"4F",  -- 79
        32566 => X"42",  -- 66
        32567 => X"3E",  -- 62
        32568 => X"3C",  -- 60
        32569 => X"45",  -- 69
        32570 => X"6B",  -- 107
        32571 => X"91",  -- 145
        32572 => X"9A",  -- 154
        32573 => X"9E",  -- 158
        32574 => X"A1",  -- 161
        32575 => X"9B",  -- 155
        32576 => X"96",  -- 150
        32577 => X"A6",  -- 166
        32578 => X"99",  -- 153
        32579 => X"9E",  -- 158
        32580 => X"A6",  -- 166
        32581 => X"B7",  -- 183
        32582 => X"AE",  -- 174
        32583 => X"B6",  -- 182
        32584 => X"AD",  -- 173
        32585 => X"AB",  -- 171
        32586 => X"B4",  -- 180
        32587 => X"AE",  -- 174
        32588 => X"A9",  -- 169
        32589 => X"99",  -- 153
        32590 => X"B3",  -- 179
        32591 => X"B5",  -- 181
        32592 => X"B5",  -- 181
        32593 => X"AC",  -- 172
        32594 => X"A8",  -- 168
        32595 => X"A5",  -- 165
        32596 => X"96",  -- 150
        32597 => X"A0",  -- 160
        32598 => X"8E",  -- 142
        32599 => X"8A",  -- 138
        32600 => X"84",  -- 132
        32601 => X"88",  -- 136
        32602 => X"83",  -- 131
        32603 => X"80",  -- 128
        32604 => X"74",  -- 116
        32605 => X"73",  -- 115
        32606 => X"89",  -- 137
        32607 => X"8E",  -- 142
        32608 => X"90",  -- 144
        32609 => X"98",  -- 152
        32610 => X"98",  -- 152
        32611 => X"8F",  -- 143
        32612 => X"91",  -- 145
        32613 => X"9D",  -- 157
        32614 => X"A7",  -- 167
        32615 => X"A6",  -- 166
        32616 => X"B4",  -- 180
        32617 => X"B4",  -- 180
        32618 => X"B8",  -- 184
        32619 => X"BD",  -- 189
        32620 => X"B7",  -- 183
        32621 => X"AB",  -- 171
        32622 => X"AB",  -- 171
        32623 => X"B4",  -- 180
        32624 => X"BC",  -- 188
        32625 => X"C3",  -- 195
        32626 => X"C7",  -- 199
        32627 => X"C3",  -- 195
        32628 => X"BD",  -- 189
        32629 => X"B9",  -- 185
        32630 => X"B7",  -- 183
        32631 => X"B4",  -- 180
        32632 => X"BD",  -- 189
        32633 => X"BD",  -- 189
        32634 => X"BC",  -- 188
        32635 => X"BD",  -- 189
        32636 => X"C1",  -- 193
        32637 => X"BC",  -- 188
        32638 => X"AE",  -- 174
        32639 => X"9F",  -- 159
        32640 => X"5B",  -- 91
        32641 => X"5B",  -- 91
        32642 => X"5A",  -- 90
        32643 => X"5B",  -- 91
        32644 => X"60",  -- 96
        32645 => X"67",  -- 103
        32646 => X"6C",  -- 108
        32647 => X"70",  -- 112
        32648 => X"6F",  -- 111
        32649 => X"69",  -- 105
        32650 => X"62",  -- 98
        32651 => X"60",  -- 96
        32652 => X"60",  -- 96
        32653 => X"5E",  -- 94
        32654 => X"5A",  -- 90
        32655 => X"55",  -- 85
        32656 => X"52",  -- 82
        32657 => X"52",  -- 82
        32658 => X"52",  -- 82
        32659 => X"52",  -- 82
        32660 => X"53",  -- 83
        32661 => X"54",  -- 84
        32662 => X"55",  -- 85
        32663 => X"56",  -- 86
        32664 => X"56",  -- 86
        32665 => X"53",  -- 83
        32666 => X"52",  -- 82
        32667 => X"56",  -- 86
        32668 => X"54",  -- 84
        32669 => X"52",  -- 82
        32670 => X"5E",  -- 94
        32671 => X"6C",  -- 108
        32672 => X"71",  -- 113
        32673 => X"6B",  -- 107
        32674 => X"53",  -- 83
        32675 => X"2F",  -- 47
        32676 => X"15",  -- 21
        32677 => X"0D",  -- 13
        32678 => X"0E",  -- 14
        32679 => X"0E",  -- 14
        32680 => X"46",  -- 70
        32681 => X"78",  -- 120
        32682 => X"50",  -- 80
        32683 => X"1F",  -- 31
        32684 => X"13",  -- 19
        32685 => X"10",  -- 16
        32686 => X"23",  -- 35
        32687 => X"26",  -- 38
        32688 => X"3A",  -- 58
        32689 => X"3F",  -- 63
        32690 => X"3F",  -- 63
        32691 => X"2D",  -- 45
        32692 => X"13",  -- 19
        32693 => X"1F",  -- 31
        32694 => X"6B",  -- 107
        32695 => X"BA",  -- 186
        32696 => X"B2",  -- 178
        32697 => X"76",  -- 118
        32698 => X"4F",  -- 79
        32699 => X"46",  -- 70
        32700 => X"42",  -- 66
        32701 => X"50",  -- 80
        32702 => X"81",  -- 129
        32703 => X"BB",  -- 187
        32704 => X"AE",  -- 174
        32705 => X"53",  -- 83
        32706 => X"3E",  -- 62
        32707 => X"80",  -- 128
        32708 => X"73",  -- 115
        32709 => X"79",  -- 121
        32710 => X"98",  -- 152
        32711 => X"AD",  -- 173
        32712 => X"D0",  -- 208
        32713 => X"C9",  -- 201
        32714 => X"C5",  -- 197
        32715 => X"C2",  -- 194
        32716 => X"9E",  -- 158
        32717 => X"68",  -- 104
        32718 => X"3F",  -- 63
        32719 => X"2A",  -- 42
        32720 => X"4D",  -- 77
        32721 => X"53",  -- 83
        32722 => X"62",  -- 98
        32723 => X"7D",  -- 125
        32724 => X"74",  -- 116
        32725 => X"77",  -- 119
        32726 => X"63",  -- 99
        32727 => X"5C",  -- 92
        32728 => X"52",  -- 82
        32729 => X"12",  -- 18
        32730 => X"2A",  -- 42
        32731 => X"69",  -- 105
        32732 => X"4A",  -- 74
        32733 => X"4E",  -- 78
        32734 => X"52",  -- 82
        32735 => X"58",  -- 88
        32736 => X"5E",  -- 94
        32737 => X"60",  -- 96
        32738 => X"42",  -- 66
        32739 => X"46",  -- 70
        32740 => X"0F",  -- 15
        32741 => X"45",  -- 69
        32742 => X"4D",  -- 77
        32743 => X"1E",  -- 30
        32744 => X"31",  -- 49
        32745 => X"65",  -- 101
        32746 => X"8C",  -- 140
        32747 => X"4A",  -- 74
        32748 => X"26",  -- 38
        32749 => X"54",  -- 84
        32750 => X"5B",  -- 91
        32751 => X"53",  -- 83
        32752 => X"90",  -- 144
        32753 => X"B4",  -- 180
        32754 => X"C5",  -- 197
        32755 => X"C8",  -- 200
        32756 => X"C5",  -- 197
        32757 => X"C2",  -- 194
        32758 => X"90",  -- 144
        32759 => X"7F",  -- 127
        32760 => X"C1",  -- 193
        32761 => X"D0",  -- 208
        32762 => X"DA",  -- 218
        32763 => X"E8",  -- 232
        32764 => X"DD",  -- 221
        32765 => X"D5",  -- 213
        32766 => X"C6",  -- 198
        32767 => X"85",  -- 133
        32768 => X"60",  -- 96
        32769 => X"8A",  -- 138
        32770 => X"BD",  -- 189
        32771 => X"D9",  -- 217
        32772 => X"CA",  -- 202
        32773 => X"E0",  -- 224
        32774 => X"DB",  -- 219
        32775 => X"C5",  -- 197
        32776 => X"7B",  -- 123
        32777 => X"32",  -- 50
        32778 => X"38",  -- 56
        32779 => X"4D",  -- 77
        32780 => X"79",  -- 121
        32781 => X"92",  -- 146
        32782 => X"9E",  -- 158
        32783 => X"B5",  -- 181
        32784 => X"BF",  -- 191
        32785 => X"B0",  -- 176
        32786 => X"97",  -- 151
        32787 => X"60",  -- 96
        32788 => X"3A",  -- 58
        32789 => X"31",  -- 49
        32790 => X"4B",  -- 75
        32791 => X"8D",  -- 141
        32792 => X"69",  -- 105
        32793 => X"1E",  -- 30
        32794 => X"0B",  -- 11
        32795 => X"0C",  -- 12
        32796 => X"1C",  -- 28
        32797 => X"2F",  -- 47
        32798 => X"63",  -- 99
        32799 => X"92",  -- 146
        32800 => X"BF",  -- 191
        32801 => X"BB",  -- 187
        32802 => X"B2",  -- 178
        32803 => X"AE",  -- 174
        32804 => X"B3",  -- 179
        32805 => X"BC",  -- 188
        32806 => X"BC",  -- 188
        32807 => X"B7",  -- 183
        32808 => X"C4",  -- 196
        32809 => X"C6",  -- 198
        32810 => X"C5",  -- 197
        32811 => X"BD",  -- 189
        32812 => X"B1",  -- 177
        32813 => X"A5",  -- 165
        32814 => X"9E",  -- 158
        32815 => X"9A",  -- 154
        32816 => X"9F",  -- 159
        32817 => X"96",  -- 150
        32818 => X"91",  -- 145
        32819 => X"93",  -- 147
        32820 => X"88",  -- 136
        32821 => X"72",  -- 114
        32822 => X"62",  -- 98
        32823 => X"5D",  -- 93
        32824 => X"4D",  -- 77
        32825 => X"34",  -- 52
        32826 => X"20",  -- 32
        32827 => X"28",  -- 40
        32828 => X"40",  -- 64
        32829 => X"59",  -- 89
        32830 => X"6E",  -- 110
        32831 => X"7D",  -- 125
        32832 => X"7E",  -- 126
        32833 => X"67",  -- 103
        32834 => X"56",  -- 86
        32835 => X"52",  -- 82
        32836 => X"4C",  -- 76
        32837 => X"44",  -- 68
        32838 => X"40",  -- 64
        32839 => X"3D",  -- 61
        32840 => X"27",  -- 39
        32841 => X"3C",  -- 60
        32842 => X"58",  -- 88
        32843 => X"6F",  -- 111
        32844 => X"84",  -- 132
        32845 => X"96",  -- 150
        32846 => X"A1",  -- 161
        32847 => X"A3",  -- 163
        32848 => X"AB",  -- 171
        32849 => X"AB",  -- 171
        32850 => X"AD",  -- 173
        32851 => X"AE",  -- 174
        32852 => X"AC",  -- 172
        32853 => X"AA",  -- 170
        32854 => X"AE",  -- 174
        32855 => X"B5",  -- 181
        32856 => X"BE",  -- 190
        32857 => X"BB",  -- 187
        32858 => X"B5",  -- 181
        32859 => X"B0",  -- 176
        32860 => X"B5",  -- 181
        32861 => X"BC",  -- 188
        32862 => X"B6",  -- 182
        32863 => X"A8",  -- 168
        32864 => X"90",  -- 144
        32865 => X"8B",  -- 139
        32866 => X"97",  -- 151
        32867 => X"A9",  -- 169
        32868 => X"AE",  -- 174
        32869 => X"B3",  -- 179
        32870 => X"BA",  -- 186
        32871 => X"BC",  -- 188
        32872 => X"BA",  -- 186
        32873 => X"BC",  -- 188
        32874 => X"BD",  -- 189
        32875 => X"BD",  -- 189
        32876 => X"BC",  -- 188
        32877 => X"BB",  -- 187
        32878 => X"BB",  -- 187
        32879 => X"BC",  -- 188
        32880 => X"BA",  -- 186
        32881 => X"A8",  -- 168
        32882 => X"94",  -- 148
        32883 => X"70",  -- 112
        32884 => X"5D",  -- 93
        32885 => X"5A",  -- 90
        32886 => X"43",  -- 67
        32887 => X"34",  -- 52
        32888 => X"45",  -- 69
        32889 => X"55",  -- 85
        32890 => X"76",  -- 118
        32891 => X"94",  -- 148
        32892 => X"9C",  -- 156
        32893 => X"97",  -- 151
        32894 => X"94",  -- 148
        32895 => X"96",  -- 150
        32896 => X"8D",  -- 141
        32897 => X"A7",  -- 167
        32898 => X"A1",  -- 161
        32899 => X"A7",  -- 167
        32900 => X"AE",  -- 174
        32901 => X"B4",  -- 180
        32902 => X"A3",  -- 163
        32903 => X"AC",  -- 172
        32904 => X"AE",  -- 174
        32905 => X"AB",  -- 171
        32906 => X"AC",  -- 172
        32907 => X"B2",  -- 178
        32908 => X"A7",  -- 167
        32909 => X"9A",  -- 154
        32910 => X"B4",  -- 180
        32911 => X"AF",  -- 175
        32912 => X"AE",  -- 174
        32913 => X"AA",  -- 170
        32914 => X"9F",  -- 159
        32915 => X"95",  -- 149
        32916 => X"8C",  -- 140
        32917 => X"9E",  -- 158
        32918 => X"8E",  -- 142
        32919 => X"85",  -- 133
        32920 => X"7F",  -- 127
        32921 => X"84",  -- 132
        32922 => X"76",  -- 118
        32923 => X"7C",  -- 124
        32924 => X"7F",  -- 127
        32925 => X"77",  -- 119
        32926 => X"87",  -- 135
        32927 => X"91",  -- 145
        32928 => X"9D",  -- 157
        32929 => X"9E",  -- 158
        32930 => X"9E",  -- 158
        32931 => X"97",  -- 151
        32932 => X"96",  -- 150
        32933 => X"9C",  -- 156
        32934 => X"A5",  -- 165
        32935 => X"AC",  -- 172
        32936 => X"BC",  -- 188
        32937 => X"BB",  -- 187
        32938 => X"BF",  -- 191
        32939 => X"BE",  -- 190
        32940 => X"AC",  -- 172
        32941 => X"99",  -- 153
        32942 => X"9E",  -- 158
        32943 => X"AE",  -- 174
        32944 => X"BD",  -- 189
        32945 => X"C5",  -- 197
        32946 => X"CA",  -- 202
        32947 => X"C9",  -- 201
        32948 => X"C3",  -- 195
        32949 => X"BF",  -- 191
        32950 => X"BB",  -- 187
        32951 => X"B6",  -- 182
        32952 => X"BA",  -- 186
        32953 => X"BC",  -- 188
        32954 => X"BF",  -- 191
        32955 => X"C1",  -- 193
        32956 => X"C1",  -- 193
        32957 => X"BC",  -- 188
        32958 => X"AF",  -- 175
        32959 => X"A0",  -- 160
        32960 => X"59",  -- 89
        32961 => X"59",  -- 89
        32962 => X"59",  -- 89
        32963 => X"5B",  -- 91
        32964 => X"61",  -- 97
        32965 => X"67",  -- 103
        32966 => X"6B",  -- 107
        32967 => X"6F",  -- 111
        32968 => X"74",  -- 116
        32969 => X"6E",  -- 110
        32970 => X"68",  -- 104
        32971 => X"66",  -- 102
        32972 => X"67",  -- 103
        32973 => X"66",  -- 102
        32974 => X"61",  -- 97
        32975 => X"5B",  -- 91
        32976 => X"53",  -- 83
        32977 => X"50",  -- 80
        32978 => X"4C",  -- 76
        32979 => X"4A",  -- 74
        32980 => X"49",  -- 73
        32981 => X"4C",  -- 76
        32982 => X"4F",  -- 79
        32983 => X"52",  -- 82
        32984 => X"52",  -- 82
        32985 => X"4F",  -- 79
        32986 => X"53",  -- 83
        32987 => X"58",  -- 88
        32988 => X"57",  -- 87
        32989 => X"58",  -- 88
        32990 => X"64",  -- 100
        32991 => X"75",  -- 117
        32992 => X"5F",  -- 95
        32993 => X"66",  -- 102
        32994 => X"53",  -- 83
        32995 => X"26",  -- 38
        32996 => X"07",  -- 7
        32997 => X"08",  -- 8
        32998 => X"0F",  -- 15
        32999 => X"0D",  -- 13
        33000 => X"50",  -- 80
        33001 => X"72",  -- 114
        33002 => X"43",  -- 67
        33003 => X"21",  -- 33
        33004 => X"18",  -- 24
        33005 => X"0D",  -- 13
        33006 => X"1E",  -- 30
        33007 => X"1D",  -- 29
        33008 => X"29",  -- 41
        33009 => X"1B",  -- 27
        33010 => X"10",  -- 16
        33011 => X"10",  -- 16
        33012 => X"1F",  -- 31
        33013 => X"48",  -- 72
        33014 => X"8B",  -- 139
        33015 => X"C4",  -- 196
        33016 => X"C3",  -- 195
        33017 => X"C0",  -- 192
        33018 => X"B2",  -- 178
        33019 => X"AF",  -- 175
        33020 => X"BF",  -- 191
        33021 => X"B0",  -- 176
        33022 => X"98",  -- 152
        33023 => X"AD",  -- 173
        33024 => X"BA",  -- 186
        33025 => X"B8",  -- 184
        33026 => X"74",  -- 116
        33027 => X"78",  -- 120
        33028 => X"7B",  -- 123
        33029 => X"66",  -- 102
        33030 => X"96",  -- 150
        33031 => X"B0",  -- 176
        33032 => X"B2",  -- 178
        33033 => X"CD",  -- 205
        33034 => X"C4",  -- 196
        33035 => X"9E",  -- 158
        33036 => X"91",  -- 145
        33037 => X"51",  -- 81
        33038 => X"0C",  -- 12
        33039 => X"2C",  -- 44
        33040 => X"7E",  -- 126
        33041 => X"66",  -- 102
        33042 => X"6A",  -- 106
        33043 => X"67",  -- 103
        33044 => X"7B",  -- 123
        33045 => X"78",  -- 120
        33046 => X"6C",  -- 108
        33047 => X"52",  -- 82
        33048 => X"27",  -- 39
        33049 => X"1F",  -- 31
        33050 => X"62",  -- 98
        33051 => X"76",  -- 118
        33052 => X"23",  -- 35
        33053 => X"4E",  -- 78
        33054 => X"66",  -- 102
        33055 => X"58",  -- 88
        33056 => X"64",  -- 100
        33057 => X"5D",  -- 93
        33058 => X"49",  -- 73
        33059 => X"3A",  -- 58
        33060 => X"1A",  -- 26
        33061 => X"38",  -- 56
        33062 => X"51",  -- 81
        33063 => X"22",  -- 34
        33064 => X"1F",  -- 31
        33065 => X"40",  -- 64
        33066 => X"82",  -- 130
        33067 => X"81",  -- 129
        33068 => X"2F",  -- 47
        33069 => X"27",  -- 39
        33070 => X"5D",  -- 93
        33071 => X"6B",  -- 107
        33072 => X"8B",  -- 139
        33073 => X"A4",  -- 164
        33074 => X"B7",  -- 183
        33075 => X"C4",  -- 196
        33076 => X"C1",  -- 193
        33077 => X"C4",  -- 196
        33078 => X"A4",  -- 164
        33079 => X"A2",  -- 162
        33080 => X"C7",  -- 199
        33081 => X"DD",  -- 221
        33082 => X"DC",  -- 220
        33083 => X"EF",  -- 239
        33084 => X"E1",  -- 225
        33085 => X"C2",  -- 194
        33086 => X"C5",  -- 197
        33087 => X"B0",  -- 176
        33088 => X"C4",  -- 196
        33089 => X"D4",  -- 212
        33090 => X"E1",  -- 225
        33091 => X"F0",  -- 240
        33092 => X"E7",  -- 231
        33093 => X"F4",  -- 244
        33094 => X"DE",  -- 222
        33095 => X"D5",  -- 213
        33096 => X"8E",  -- 142
        33097 => X"48",  -- 72
        33098 => X"40",  -- 64
        33099 => X"2A",  -- 42
        33100 => X"2F",  -- 47
        33101 => X"44",  -- 68
        33102 => X"65",  -- 101
        33103 => X"8F",  -- 143
        33104 => X"A6",  -- 166
        33105 => X"8B",  -- 139
        33106 => X"6B",  -- 107
        33107 => X"3A",  -- 58
        33108 => X"28",  -- 40
        33109 => X"31",  -- 49
        33110 => X"54",  -- 84
        33111 => X"99",  -- 153
        33112 => X"98",  -- 152
        33113 => X"3E",  -- 62
        33114 => X"15",  -- 21
        33115 => X"09",  -- 9
        33116 => X"19",  -- 25
        33117 => X"2C",  -- 44
        33118 => X"55",  -- 85
        33119 => X"77",  -- 119
        33120 => X"AD",  -- 173
        33121 => X"BB",  -- 187
        33122 => X"B8",  -- 184
        33123 => X"A3",  -- 163
        33124 => X"9F",  -- 159
        33125 => X"B1",  -- 177
        33126 => X"BF",  -- 191
        33127 => X"BF",  -- 191
        33128 => X"C4",  -- 196
        33129 => X"C4",  -- 196
        33130 => X"C0",  -- 192
        33131 => X"BB",  -- 187
        33132 => X"B4",  -- 180
        33133 => X"AA",  -- 170
        33134 => X"A4",  -- 164
        33135 => X"9F",  -- 159
        33136 => X"A2",  -- 162
        33137 => X"A6",  -- 166
        33138 => X"98",  -- 152
        33139 => X"81",  -- 129
        33140 => X"82",  -- 130
        33141 => X"88",  -- 136
        33142 => X"6F",  -- 111
        33143 => X"47",  -- 71
        33144 => X"41",  -- 65
        33145 => X"28",  -- 40
        33146 => X"1B",  -- 27
        33147 => X"2F",  -- 47
        33148 => X"4C",  -- 76
        33149 => X"5C",  -- 92
        33150 => X"68",  -- 104
        33151 => X"71",  -- 113
        33152 => X"70",  -- 112
        33153 => X"6E",  -- 110
        33154 => X"5B",  -- 91
        33155 => X"52",  -- 82
        33156 => X"54",  -- 84
        33157 => X"3D",  -- 61
        33158 => X"29",  -- 41
        33159 => X"33",  -- 51
        33160 => X"24",  -- 36
        33161 => X"3B",  -- 59
        33162 => X"5B",  -- 91
        33163 => X"75",  -- 117
        33164 => X"8C",  -- 140
        33165 => X"A0",  -- 160
        33166 => X"AD",  -- 173
        33167 => X"B1",  -- 177
        33168 => X"A7",  -- 167
        33169 => X"A6",  -- 166
        33170 => X"AC",  -- 172
        33171 => X"B4",  -- 180
        33172 => X"B5",  -- 181
        33173 => X"AC",  -- 172
        33174 => X"A9",  -- 169
        33175 => X"AC",  -- 172
        33176 => X"B4",  -- 180
        33177 => X"B4",  -- 180
        33178 => X"B1",  -- 177
        33179 => X"AD",  -- 173
        33180 => X"B2",  -- 178
        33181 => X"B7",  -- 183
        33182 => X"AD",  -- 173
        33183 => X"9D",  -- 157
        33184 => X"A0",  -- 160
        33185 => X"98",  -- 152
        33186 => X"9F",  -- 159
        33187 => X"AA",  -- 170
        33188 => X"AC",  -- 172
        33189 => X"B2",  -- 178
        33190 => X"BC",  -- 188
        33191 => X"C2",  -- 194
        33192 => X"C0",  -- 192
        33193 => X"C1",  -- 193
        33194 => X"C2",  -- 194
        33195 => X"C1",  -- 193
        33196 => X"BE",  -- 190
        33197 => X"BA",  -- 186
        33198 => X"B8",  -- 184
        33199 => X"B7",  -- 183
        33200 => X"B1",  -- 177
        33201 => X"9B",  -- 155
        33202 => X"8D",  -- 141
        33203 => X"6F",  -- 111
        33204 => X"4C",  -- 76
        33205 => X"35",  -- 53
        33206 => X"31",  -- 49
        33207 => X"47",  -- 71
        33208 => X"51",  -- 81
        33209 => X"63",  -- 99
        33210 => X"7A",  -- 122
        33211 => X"8B",  -- 139
        33212 => X"90",  -- 144
        33213 => X"86",  -- 134
        33214 => X"82",  -- 130
        33215 => X"8E",  -- 142
        33216 => X"9C",  -- 156
        33217 => X"A1",  -- 161
        33218 => X"90",  -- 144
        33219 => X"A0",  -- 160
        33220 => X"AC",  -- 172
        33221 => X"A6",  -- 166
        33222 => X"95",  -- 149
        33223 => X"AE",  -- 174
        33224 => X"AE",  -- 174
        33225 => X"A7",  -- 167
        33226 => X"9F",  -- 159
        33227 => X"A9",  -- 169
        33228 => X"A2",  -- 162
        33229 => X"9D",  -- 157
        33230 => X"AC",  -- 172
        33231 => X"9B",  -- 155
        33232 => X"A7",  -- 167
        33233 => X"A3",  -- 163
        33234 => X"96",  -- 150
        33235 => X"89",  -- 137
        33236 => X"86",  -- 134
        33237 => X"A0",  -- 160
        33238 => X"92",  -- 146
        33239 => X"8B",  -- 139
        33240 => X"77",  -- 119
        33241 => X"7B",  -- 123
        33242 => X"67",  -- 103
        33243 => X"79",  -- 121
        33244 => X"8A",  -- 138
        33245 => X"7F",  -- 127
        33246 => X"87",  -- 135
        33247 => X"91",  -- 145
        33248 => X"9D",  -- 157
        33249 => X"9A",  -- 154
        33250 => X"9A",  -- 154
        33251 => X"9D",  -- 157
        33252 => X"9A",  -- 154
        33253 => X"99",  -- 153
        33254 => X"A6",  -- 166
        33255 => X"B7",  -- 183
        33256 => X"B8",  -- 184
        33257 => X"B8",  -- 184
        33258 => X"BC",  -- 188
        33259 => X"BA",  -- 186
        33260 => X"A4",  -- 164
        33261 => X"90",  -- 144
        33262 => X"97",  -- 151
        33263 => X"AF",  -- 175
        33264 => X"BC",  -- 188
        33265 => X"C5",  -- 197
        33266 => X"CB",  -- 203
        33267 => X"CB",  -- 203
        33268 => X"C8",  -- 200
        33269 => X"C6",  -- 198
        33270 => X"C1",  -- 193
        33271 => X"BD",  -- 189
        33272 => X"AE",  -- 174
        33273 => X"B5",  -- 181
        33274 => X"BD",  -- 189
        33275 => X"BF",  -- 191
        33276 => X"BE",  -- 190
        33277 => X"B8",  -- 184
        33278 => X"AE",  -- 174
        33279 => X"A3",  -- 163
        33280 => X"57",  -- 87
        33281 => X"5A",  -- 90
        33282 => X"5D",  -- 93
        33283 => X"5D",  -- 93
        33284 => X"5D",  -- 93
        33285 => X"5E",  -- 94
        33286 => X"5F",  -- 95
        33287 => X"62",  -- 98
        33288 => X"67",  -- 103
        33289 => X"63",  -- 99
        33290 => X"62",  -- 98
        33291 => X"68",  -- 104
        33292 => X"70",  -- 112
        33293 => X"72",  -- 114
        33294 => X"6D",  -- 109
        33295 => X"66",  -- 102
        33296 => X"5A",  -- 90
        33297 => X"53",  -- 83
        33298 => X"4B",  -- 75
        33299 => X"46",  -- 70
        33300 => X"47",  -- 71
        33301 => X"4A",  -- 74
        33302 => X"4A",  -- 74
        33303 => X"49",  -- 73
        33304 => X"49",  -- 73
        33305 => X"4F",  -- 79
        33306 => X"54",  -- 84
        33307 => X"54",  -- 84
        33308 => X"59",  -- 89
        33309 => X"61",  -- 97
        33310 => X"60",  -- 96
        33311 => X"5A",  -- 90
        33312 => X"6F",  -- 111
        33313 => X"61",  -- 97
        33314 => X"3D",  -- 61
        33315 => X"14",  -- 20
        33316 => X"0E",  -- 14
        33317 => X"0B",  -- 11
        33318 => X"08",  -- 8
        33319 => X"29",  -- 41
        33320 => X"69",  -- 105
        33321 => X"7B",  -- 123
        33322 => X"54",  -- 84
        33323 => X"1E",  -- 30
        33324 => X"12",  -- 18
        33325 => X"0E",  -- 14
        33326 => X"13",  -- 19
        33327 => X"2E",  -- 46
        33328 => X"42",  -- 66
        33329 => X"19",  -- 25
        33330 => X"0A",  -- 10
        33331 => X"16",  -- 22
        33332 => X"0F",  -- 15
        33333 => X"35",  -- 53
        33334 => X"92",  -- 146
        33335 => X"C4",  -- 196
        33336 => X"BE",  -- 190
        33337 => X"C2",  -- 194
        33338 => X"C4",  -- 196
        33339 => X"C5",  -- 197
        33340 => X"CA",  -- 202
        33341 => X"C9",  -- 201
        33342 => X"B4",  -- 180
        33343 => X"9C",  -- 156
        33344 => X"AB",  -- 171
        33345 => X"B8",  -- 184
        33346 => X"B9",  -- 185
        33347 => X"AE",  -- 174
        33348 => X"89",  -- 137
        33349 => X"57",  -- 87
        33350 => X"6E",  -- 110
        33351 => X"BF",  -- 191
        33352 => X"B7",  -- 183
        33353 => X"B9",  -- 185
        33354 => X"AC",  -- 172
        33355 => X"9F",  -- 159
        33356 => X"7D",  -- 125
        33357 => X"2E",  -- 46
        33358 => X"11",  -- 17
        33359 => X"3C",  -- 60
        33360 => X"75",  -- 117
        33361 => X"73",  -- 115
        33362 => X"54",  -- 84
        33363 => X"57",  -- 87
        33364 => X"69",  -- 105
        33365 => X"71",  -- 113
        33366 => X"61",  -- 97
        33367 => X"2A",  -- 42
        33368 => X"23",  -- 35
        33369 => X"4F",  -- 79
        33370 => X"72",  -- 114
        33371 => X"4A",  -- 74
        33372 => X"29",  -- 41
        33373 => X"5B",  -- 91
        33374 => X"5C",  -- 92
        33375 => X"62",  -- 98
        33376 => X"5A",  -- 90
        33377 => X"69",  -- 105
        33378 => X"2F",  -- 47
        33379 => X"31",  -- 49
        33380 => X"35",  -- 53
        33381 => X"1F",  -- 31
        33382 => X"62",  -- 98
        33383 => X"2A",  -- 42
        33384 => X"1E",  -- 30
        33385 => X"4E",  -- 78
        33386 => X"79",  -- 121
        33387 => X"88",  -- 136
        33388 => X"44",  -- 68
        33389 => X"0B",  -- 11
        33390 => X"33",  -- 51
        33391 => X"79",  -- 121
        33392 => X"81",  -- 129
        33393 => X"9F",  -- 159
        33394 => X"B8",  -- 184
        33395 => X"C2",  -- 194
        33396 => X"CA",  -- 202
        33397 => X"C9",  -- 201
        33398 => X"B8",  -- 184
        33399 => X"A2",  -- 162
        33400 => X"D3",  -- 211
        33401 => X"DB",  -- 219
        33402 => X"DC",  -- 220
        33403 => X"E4",  -- 228
        33404 => X"CE",  -- 206
        33405 => X"C2",  -- 194
        33406 => X"D9",  -- 217
        33407 => X"D1",  -- 209
        33408 => X"DC",  -- 220
        33409 => X"EE",  -- 238
        33410 => X"EB",  -- 235
        33411 => X"E8",  -- 232
        33412 => X"EB",  -- 235
        33413 => X"ED",  -- 237
        33414 => X"E9",  -- 233
        33415 => X"CE",  -- 206
        33416 => X"7A",  -- 122
        33417 => X"58",  -- 88
        33418 => X"3A",  -- 58
        33419 => X"18",  -- 24
        33420 => X"1A",  -- 26
        33421 => X"28",  -- 40
        33422 => X"37",  -- 55
        33423 => X"66",  -- 102
        33424 => X"8D",  -- 141
        33425 => X"78",  -- 120
        33426 => X"4C",  -- 76
        33427 => X"26",  -- 38
        33428 => X"27",  -- 39
        33429 => X"34",  -- 52
        33430 => X"52",  -- 82
        33431 => X"8D",  -- 141
        33432 => X"84",  -- 132
        33433 => X"3B",  -- 59
        33434 => X"12",  -- 18
        33435 => X"11",  -- 17
        33436 => X"0F",  -- 15
        33437 => X"20",  -- 32
        33438 => X"4E",  -- 78
        33439 => X"6F",  -- 111
        33440 => X"A0",  -- 160
        33441 => X"B7",  -- 183
        33442 => X"BC",  -- 188
        33443 => X"AF",  -- 175
        33444 => X"AB",  -- 171
        33445 => X"B3",  -- 179
        33446 => X"BC",  -- 188
        33447 => X"C6",  -- 198
        33448 => X"C6",  -- 198
        33449 => X"CB",  -- 203
        33450 => X"C8",  -- 200
        33451 => X"BA",  -- 186
        33452 => X"B0",  -- 176
        33453 => X"AD",  -- 173
        33454 => X"AC",  -- 172
        33455 => X"AA",  -- 170
        33456 => X"9B",  -- 155
        33457 => X"A3",  -- 163
        33458 => X"A5",  -- 165
        33459 => X"90",  -- 144
        33460 => X"73",  -- 115
        33461 => X"6C",  -- 108
        33462 => X"6D",  -- 109
        33463 => X"67",  -- 103
        33464 => X"3C",  -- 60
        33465 => X"20",  -- 32
        33466 => X"18",  -- 24
        33467 => X"2E",  -- 46
        33468 => X"48",  -- 72
        33469 => X"5C",  -- 92
        33470 => X"6A",  -- 106
        33471 => X"6E",  -- 110
        33472 => X"6D",  -- 109
        33473 => X"64",  -- 100
        33474 => X"5A",  -- 90
        33475 => X"51",  -- 81
        33476 => X"46",  -- 70
        33477 => X"35",  -- 53
        33478 => X"25",  -- 37
        33479 => X"1D",  -- 29
        33480 => X"20",  -- 32
        33481 => X"27",  -- 39
        33482 => X"50",  -- 80
        33483 => X"7B",  -- 123
        33484 => X"8B",  -- 139
        33485 => X"99",  -- 153
        33486 => X"AD",  -- 173
        33487 => X"B5",  -- 181
        33488 => X"B0",  -- 176
        33489 => X"AE",  -- 174
        33490 => X"B3",  -- 179
        33491 => X"B8",  -- 184
        33492 => X"B6",  -- 182
        33493 => X"AE",  -- 174
        33494 => X"AF",  -- 175
        33495 => X"B6",  -- 182
        33496 => X"B9",  -- 185
        33497 => X"BA",  -- 186
        33498 => X"B5",  -- 181
        33499 => X"AA",  -- 170
        33500 => X"AA",  -- 170
        33501 => X"B0",  -- 176
        33502 => X"B1",  -- 177
        33503 => X"AB",  -- 171
        33504 => X"93",  -- 147
        33505 => X"9C",  -- 156
        33506 => X"A7",  -- 167
        33507 => X"B0",  -- 176
        33508 => X"B3",  -- 179
        33509 => X"B4",  -- 180
        33510 => X"B4",  -- 180
        33511 => X"B6",  -- 182
        33512 => X"B5",  -- 181
        33513 => X"BA",  -- 186
        33514 => X"BD",  -- 189
        33515 => X"BA",  -- 186
        33516 => X"B7",  -- 183
        33517 => X"B6",  -- 182
        33518 => X"B5",  -- 181
        33519 => X"B1",  -- 177
        33520 => X"B7",  -- 183
        33521 => X"9C",  -- 156
        33522 => X"87",  -- 135
        33523 => X"78",  -- 120
        33524 => X"5E",  -- 94
        33525 => X"3B",  -- 59
        33526 => X"30",  -- 48
        33527 => X"39",  -- 57
        33528 => X"57",  -- 87
        33529 => X"67",  -- 103
        33530 => X"6B",  -- 107
        33531 => X"75",  -- 117
        33532 => X"79",  -- 121
        33533 => X"7A",  -- 122
        33534 => X"82",  -- 130
        33535 => X"7C",  -- 124
        33536 => X"9C",  -- 156
        33537 => X"9C",  -- 156
        33538 => X"91",  -- 145
        33539 => X"9A",  -- 154
        33540 => X"AD",  -- 173
        33541 => X"A1",  -- 161
        33542 => X"91",  -- 145
        33543 => X"A1",  -- 161
        33544 => X"AA",  -- 170
        33545 => X"91",  -- 145
        33546 => X"A3",  -- 163
        33547 => X"AE",  -- 174
        33548 => X"8E",  -- 142
        33549 => X"9E",  -- 158
        33550 => X"97",  -- 151
        33551 => X"96",  -- 150
        33552 => X"9A",  -- 154
        33553 => X"A2",  -- 162
        33554 => X"8C",  -- 140
        33555 => X"8B",  -- 139
        33556 => X"8B",  -- 139
        33557 => X"86",  -- 134
        33558 => X"8C",  -- 140
        33559 => X"89",  -- 137
        33560 => X"69",  -- 105
        33561 => X"73",  -- 115
        33562 => X"77",  -- 119
        33563 => X"75",  -- 117
        33564 => X"7E",  -- 126
        33565 => X"92",  -- 146
        33566 => X"98",  -- 152
        33567 => X"91",  -- 145
        33568 => X"95",  -- 149
        33569 => X"9B",  -- 155
        33570 => X"9E",  -- 158
        33571 => X"A2",  -- 162
        33572 => X"A9",  -- 169
        33573 => X"AC",  -- 172
        33574 => X"AA",  -- 170
        33575 => X"A2",  -- 162
        33576 => X"B2",  -- 178
        33577 => X"BE",  -- 190
        33578 => X"B3",  -- 179
        33579 => X"A1",  -- 161
        33580 => X"9D",  -- 157
        33581 => X"98",  -- 152
        33582 => X"9B",  -- 155
        33583 => X"AB",  -- 171
        33584 => X"BA",  -- 186
        33585 => X"C2",  -- 194
        33586 => X"C9",  -- 201
        33587 => X"CD",  -- 205
        33588 => X"CE",  -- 206
        33589 => X"CD",  -- 205
        33590 => X"C6",  -- 198
        33591 => X"C1",  -- 193
        33592 => X"B6",  -- 182
        33593 => X"B7",  -- 183
        33594 => X"B9",  -- 185
        33595 => X"B9",  -- 185
        33596 => X"B7",  -- 183
        33597 => X"B3",  -- 179
        33598 => X"A7",  -- 167
        33599 => X"9E",  -- 158
        33600 => X"56",  -- 86
        33601 => X"59",  -- 89
        33602 => X"5C",  -- 92
        33603 => X"5C",  -- 92
        33604 => X"5C",  -- 92
        33605 => X"5B",  -- 91
        33606 => X"5C",  -- 92
        33607 => X"5F",  -- 95
        33608 => X"5E",  -- 94
        33609 => X"5B",  -- 91
        33610 => X"5B",  -- 91
        33611 => X"62",  -- 98
        33612 => X"6D",  -- 109
        33613 => X"72",  -- 114
        33614 => X"70",  -- 112
        33615 => X"6B",  -- 107
        33616 => X"62",  -- 98
        33617 => X"5B",  -- 91
        33618 => X"51",  -- 81
        33619 => X"4B",  -- 75
        33620 => X"4B",  -- 75
        33621 => X"4C",  -- 76
        33622 => X"4B",  -- 75
        33623 => X"4A",  -- 74
        33624 => X"4C",  -- 76
        33625 => X"4F",  -- 79
        33626 => X"50",  -- 80
        33627 => X"53",  -- 83
        33628 => X"5C",  -- 92
        33629 => X"63",  -- 99
        33630 => X"61",  -- 97
        33631 => X"5E",  -- 94
        33632 => X"64",  -- 100
        33633 => X"4F",  -- 79
        33634 => X"2D",  -- 45
        33635 => X"0E",  -- 14
        33636 => X"0B",  -- 11
        33637 => X"04",  -- 4
        33638 => X"07",  -- 7
        33639 => X"36",  -- 54
        33640 => X"71",  -- 113
        33641 => X"7B",  -- 123
        33642 => X"51",  -- 81
        33643 => X"1B",  -- 27
        33644 => X"11",  -- 17
        33645 => X"0E",  -- 14
        33646 => X"1A",  -- 26
        33647 => X"40",  -- 64
        33648 => X"59",  -- 89
        33649 => X"2F",  -- 47
        33650 => X"13",  -- 19
        33651 => X"13",  -- 19
        33652 => X"0B",  -- 11
        33653 => X"2A",  -- 42
        33654 => X"7F",  -- 127
        33655 => X"B5",  -- 181
        33656 => X"B9",  -- 185
        33657 => X"BC",  -- 188
        33658 => X"BC",  -- 188
        33659 => X"BE",  -- 190
        33660 => X"C7",  -- 199
        33661 => X"CA",  -- 202
        33662 => X"BD",  -- 189
        33663 => X"AB",  -- 171
        33664 => X"B5",  -- 181
        33665 => X"B6",  -- 182
        33666 => X"B1",  -- 177
        33667 => X"B0",  -- 176
        33668 => X"9C",  -- 156
        33669 => X"6A",  -- 106
        33670 => X"5C",  -- 92
        33671 => X"81",  -- 129
        33672 => X"A5",  -- 165
        33673 => X"A6",  -- 166
        33674 => X"95",  -- 149
        33675 => X"82",  -- 130
        33676 => X"63",  -- 99
        33677 => X"21",  -- 33
        33678 => X"0D",  -- 13
        33679 => X"36",  -- 54
        33680 => X"47",  -- 71
        33681 => X"69",  -- 105
        33682 => X"6C",  -- 108
        33683 => X"5F",  -- 95
        33684 => X"6C",  -- 108
        33685 => X"60",  -- 96
        33686 => X"35",  -- 53
        33687 => X"26",  -- 38
        33688 => X"3D",  -- 61
        33689 => X"53",  -- 83
        33690 => X"70",  -- 112
        33691 => X"55",  -- 85
        33692 => X"48",  -- 72
        33693 => X"6E",  -- 110
        33694 => X"63",  -- 99
        33695 => X"59",  -- 89
        33696 => X"4D",  -- 77
        33697 => X"6D",  -- 109
        33698 => X"46",  -- 70
        33699 => X"1B",  -- 27
        33700 => X"23",  -- 35
        33701 => X"47",  -- 71
        33702 => X"54",  -- 84
        33703 => X"4A",  -- 74
        33704 => X"3C",  -- 60
        33705 => X"63",  -- 99
        33706 => X"7F",  -- 127
        33707 => X"8B",  -- 139
        33708 => X"50",  -- 80
        33709 => X"0C",  -- 12
        33710 => X"1B",  -- 27
        33711 => X"51",  -- 81
        33712 => X"83",  -- 131
        33713 => X"91",  -- 145
        33714 => X"A6",  -- 166
        33715 => X"BB",  -- 187
        33716 => X"C2",  -- 194
        33717 => X"A2",  -- 162
        33718 => X"80",  -- 128
        33719 => X"8D",  -- 141
        33720 => X"C0",  -- 192
        33721 => X"D1",  -- 209
        33722 => X"CE",  -- 206
        33723 => X"C1",  -- 193
        33724 => X"B5",  -- 181
        33725 => X"C0",  -- 192
        33726 => X"D5",  -- 213
        33727 => X"D0",  -- 208
        33728 => X"DA",  -- 218
        33729 => X"DC",  -- 220
        33730 => X"D6",  -- 214
        33731 => X"EC",  -- 236
        33732 => X"FB",  -- 251
        33733 => X"E8",  -- 232
        33734 => X"DC",  -- 220
        33735 => X"D6",  -- 214
        33736 => X"8B",  -- 139
        33737 => X"42",  -- 66
        33738 => X"23",  -- 35
        33739 => X"19",  -- 25
        33740 => X"0C",  -- 12
        33741 => X"22",  -- 34
        33742 => X"4E",  -- 78
        33743 => X"6E",  -- 110
        33744 => X"79",  -- 121
        33745 => X"54",  -- 84
        33746 => X"2C",  -- 44
        33747 => X"1C",  -- 28
        33748 => X"2D",  -- 45
        33749 => X"42",  -- 66
        33750 => X"61",  -- 97
        33751 => X"8B",  -- 139
        33752 => X"95",  -- 149
        33753 => X"58",  -- 88
        33754 => X"1D",  -- 29
        33755 => X"0B",  -- 11
        33756 => X"0F",  -- 15
        33757 => X"14",  -- 20
        33758 => X"37",  -- 55
        33759 => X"68",  -- 104
        33760 => X"8E",  -- 142
        33761 => X"AA",  -- 170
        33762 => X"B7",  -- 183
        33763 => X"AF",  -- 175
        33764 => X"B2",  -- 178
        33765 => X"BA",  -- 186
        33766 => X"BD",  -- 189
        33767 => X"BD",  -- 189
        33768 => X"CA",  -- 202
        33769 => X"C9",  -- 201
        33770 => X"C2",  -- 194
        33771 => X"BB",  -- 187
        33772 => X"BB",  -- 187
        33773 => X"BA",  -- 186
        33774 => X"B1",  -- 177
        33775 => X"A3",  -- 163
        33776 => X"A3",  -- 163
        33777 => X"98",  -- 152
        33778 => X"94",  -- 148
        33779 => X"8E",  -- 142
        33780 => X"77",  -- 119
        33781 => X"61",  -- 97
        33782 => X"5D",  -- 93
        33783 => X"5C",  -- 92
        33784 => X"4F",  -- 79
        33785 => X"2B",  -- 43
        33786 => X"16",  -- 22
        33787 => X"24",  -- 36
        33788 => X"42",  -- 66
        33789 => X"5F",  -- 95
        33790 => X"6F",  -- 111
        33791 => X"6D",  -- 109
        33792 => X"6E",  -- 110
        33793 => X"5F",  -- 95
        33794 => X"4C",  -- 76
        33795 => X"3F",  -- 63
        33796 => X"3B",  -- 59
        33797 => X"33",  -- 51
        33798 => X"25",  -- 37
        33799 => X"19",  -- 25
        33800 => X"2A",  -- 42
        33801 => X"37",  -- 55
        33802 => X"58",  -- 88
        33803 => X"7B",  -- 123
        33804 => X"90",  -- 144
        33805 => X"9D",  -- 157
        33806 => X"AA",  -- 170
        33807 => X"AE",  -- 174
        33808 => X"B4",  -- 180
        33809 => X"AB",  -- 171
        33810 => X"A7",  -- 167
        33811 => X"AE",  -- 174
        33812 => X"B7",  -- 183
        33813 => X"B8",  -- 184
        33814 => X"B2",  -- 178
        33815 => X"AD",  -- 173
        33816 => X"A4",  -- 164
        33817 => X"B3",  -- 179
        33818 => X"BF",  -- 191
        33819 => X"BD",  -- 189
        33820 => X"BA",  -- 186
        33821 => X"B8",  -- 184
        33822 => X"B3",  -- 179
        33823 => X"AB",  -- 171
        33824 => X"9C",  -- 156
        33825 => X"A1",  -- 161
        33826 => X"A8",  -- 168
        33827 => X"AA",  -- 170
        33828 => X"AB",  -- 171
        33829 => X"AC",  -- 172
        33830 => X"AE",  -- 174
        33831 => X"AF",  -- 175
        33832 => X"AD",  -- 173
        33833 => X"AF",  -- 175
        33834 => X"AF",  -- 175
        33835 => X"AB",  -- 171
        33836 => X"AA",  -- 170
        33837 => X"AA",  -- 170
        33838 => X"A8",  -- 168
        33839 => X"A3",  -- 163
        33840 => X"9F",  -- 159
        33841 => X"8C",  -- 140
        33842 => X"75",  -- 117
        33843 => X"5E",  -- 94
        33844 => X"49",  -- 73
        33845 => X"3B",  -- 59
        33846 => X"44",  -- 68
        33847 => X"54",  -- 84
        33848 => X"5F",  -- 95
        33849 => X"6F",  -- 111
        33850 => X"6A",  -- 106
        33851 => X"63",  -- 99
        33852 => X"62",  -- 98
        33853 => X"69",  -- 105
        33854 => X"77",  -- 119
        33855 => X"6F",  -- 111
        33856 => X"8C",  -- 140
        33857 => X"98",  -- 152
        33858 => X"93",  -- 147
        33859 => X"90",  -- 144
        33860 => X"99",  -- 153
        33861 => X"8F",  -- 143
        33862 => X"84",  -- 132
        33863 => X"93",  -- 147
        33864 => X"A5",  -- 165
        33865 => X"91",  -- 145
        33866 => X"9C",  -- 156
        33867 => X"A3",  -- 163
        33868 => X"8B",  -- 139
        33869 => X"92",  -- 146
        33870 => X"86",  -- 134
        33871 => X"86",  -- 134
        33872 => X"8D",  -- 141
        33873 => X"9A",  -- 154
        33874 => X"8F",  -- 143
        33875 => X"89",  -- 137
        33876 => X"8C",  -- 140
        33877 => X"7E",  -- 126
        33878 => X"85",  -- 133
        33879 => X"7F",  -- 127
        33880 => X"6B",  -- 107
        33881 => X"6F",  -- 111
        33882 => X"76",  -- 118
        33883 => X"7E",  -- 126
        33884 => X"87",  -- 135
        33885 => X"91",  -- 145
        33886 => X"99",  -- 153
        33887 => X"9E",  -- 158
        33888 => X"9A",  -- 154
        33889 => X"9F",  -- 159
        33890 => X"A0",  -- 160
        33891 => X"A1",  -- 161
        33892 => X"A5",  -- 165
        33893 => X"AB",  -- 171
        33894 => X"AE",  -- 174
        33895 => X"AE",  -- 174
        33896 => X"B0",  -- 176
        33897 => X"C0",  -- 192
        33898 => X"B6",  -- 182
        33899 => X"97",  -- 151
        33900 => X"89",  -- 137
        33901 => X"96",  -- 150
        33902 => X"A7",  -- 167
        33903 => X"B2",  -- 178
        33904 => X"BA",  -- 186
        33905 => X"C1",  -- 193
        33906 => X"C8",  -- 200
        33907 => X"CB",  -- 203
        33908 => X"D0",  -- 208
        33909 => X"D1",  -- 209
        33910 => X"CC",  -- 204
        33911 => X"C6",  -- 198
        33912 => X"C0",  -- 192
        33913 => X"BE",  -- 190
        33914 => X"BC",  -- 188
        33915 => X"BB",  -- 187
        33916 => X"B7",  -- 183
        33917 => X"AD",  -- 173
        33918 => X"A0",  -- 160
        33919 => X"94",  -- 148
        33920 => X"54",  -- 84
        33921 => X"57",  -- 87
        33922 => X"5A",  -- 90
        33923 => X"5B",  -- 91
        33924 => X"5B",  -- 91
        33925 => X"5B",  -- 91
        33926 => X"5C",  -- 92
        33927 => X"5E",  -- 94
        33928 => X"5B",  -- 91
        33929 => X"58",  -- 88
        33930 => X"58",  -- 88
        33931 => X"5D",  -- 93
        33932 => X"66",  -- 102
        33933 => X"6B",  -- 107
        33934 => X"6A",  -- 106
        33935 => X"67",  -- 103
        33936 => X"63",  -- 99
        33937 => X"5C",  -- 92
        33938 => X"53",  -- 83
        33939 => X"4E",  -- 78
        33940 => X"4E",  -- 78
        33941 => X"4F",  -- 79
        33942 => X"4F",  -- 79
        33943 => X"4F",  -- 79
        33944 => X"4F",  -- 79
        33945 => X"4B",  -- 75
        33946 => X"4D",  -- 77
        33947 => X"57",  -- 87
        33948 => X"62",  -- 98
        33949 => X"67",  -- 103
        33950 => X"66",  -- 102
        33951 => X"66",  -- 102
        33952 => X"5C",  -- 92
        33953 => X"44",  -- 68
        33954 => X"25",  -- 37
        33955 => X"0E",  -- 14
        33956 => X"0D",  -- 13
        33957 => X"06",  -- 6
        33958 => X"12",  -- 18
        33959 => X"4F",  -- 79
        33960 => X"7C",  -- 124
        33961 => X"80",  -- 128
        33962 => X"52",  -- 82
        33963 => X"20",  -- 32
        33964 => X"10",  -- 16
        33965 => X"09",  -- 9
        33966 => X"1D",  -- 29
        33967 => X"50",  -- 80
        33968 => X"77",  -- 119
        33969 => X"4D",  -- 77
        33970 => X"1B",  -- 27
        33971 => X"0A",  -- 10
        33972 => X"05",  -- 5
        33973 => X"1A",  -- 26
        33974 => X"5F",  -- 95
        33975 => X"95",  -- 149
        33976 => X"AB",  -- 171
        33977 => X"BA",  -- 186
        33978 => X"C5",  -- 197
        33979 => X"C4",  -- 196
        33980 => X"BE",  -- 190
        33981 => X"BC",  -- 188
        33982 => X"BB",  -- 187
        33983 => X"BA",  -- 186
        33984 => X"B0",  -- 176
        33985 => X"B3",  -- 179
        33986 => X"B2",  -- 178
        33987 => X"B1",  -- 177
        33988 => X"A3",  -- 163
        33989 => X"75",  -- 117
        33990 => X"55",  -- 85
        33991 => X"5F",  -- 95
        33992 => X"85",  -- 133
        33993 => X"8C",  -- 140
        33994 => X"7D",  -- 125
        33995 => X"68",  -- 104
        33996 => X"4E",  -- 78
        33997 => X"1C",  -- 28
        33998 => X"0A",  -- 10
        33999 => X"22",  -- 34
        34000 => X"1E",  -- 30
        34001 => X"62",  -- 98
        34002 => X"81",  -- 129
        34003 => X"63",  -- 99
        34004 => X"63",  -- 99
        34005 => X"47",  -- 71
        34006 => X"11",  -- 17
        34007 => X"27",  -- 39
        34008 => X"38",  -- 56
        34009 => X"43",  -- 67
        34010 => X"66",  -- 102
        34011 => X"59",  -- 89
        34012 => X"61",  -- 97
        34013 => X"73",  -- 115
        34014 => X"61",  -- 97
        34015 => X"48",  -- 72
        34016 => X"4C",  -- 76
        34017 => X"6D",  -- 109
        34018 => X"58",  -- 88
        34019 => X"2A",  -- 42
        34020 => X"18",  -- 24
        34021 => X"49",  -- 73
        34022 => X"4F",  -- 79
        34023 => X"61",  -- 97
        34024 => X"4F",  -- 79
        34025 => X"66",  -- 102
        34026 => X"74",  -- 116
        34027 => X"7C",  -- 124
        34028 => X"5B",  -- 91
        34029 => X"10",  -- 16
        34030 => X"0F",  -- 15
        34031 => X"3D",  -- 61
        34032 => X"69",  -- 105
        34033 => X"79",  -- 121
        34034 => X"9B",  -- 155
        34035 => X"A9",  -- 169
        34036 => X"A5",  -- 165
        34037 => X"7D",  -- 125
        34038 => X"69",  -- 105
        34039 => X"A1",  -- 161
        34040 => X"C9",  -- 201
        34041 => X"D0",  -- 208
        34042 => X"CB",  -- 203
        34043 => X"AC",  -- 172
        34044 => X"A2",  -- 162
        34045 => X"A8",  -- 168
        34046 => X"A3",  -- 163
        34047 => X"A4",  -- 164
        34048 => X"A5",  -- 165
        34049 => X"CD",  -- 205
        34050 => X"E0",  -- 224
        34051 => X"D8",  -- 216
        34052 => X"D3",  -- 211
        34053 => X"E6",  -- 230
        34054 => X"DF",  -- 223
        34055 => X"9E",  -- 158
        34056 => X"5B",  -- 91
        34057 => X"2A",  -- 42
        34058 => X"12",  -- 18
        34059 => X"19",  -- 25
        34060 => X"0C",  -- 12
        34061 => X"19",  -- 25
        34062 => X"5D",  -- 93
        34063 => X"8E",  -- 142
        34064 => X"9A",  -- 154
        34065 => X"5C",  -- 92
        34066 => X"24",  -- 36
        34067 => X"18",  -- 24
        34068 => X"25",  -- 37
        34069 => X"42",  -- 66
        34070 => X"74",  -- 116
        34071 => X"9C",  -- 156
        34072 => X"9A",  -- 154
        34073 => X"65",  -- 101
        34074 => X"22",  -- 34
        34075 => X"0D",  -- 13
        34076 => X"19",  -- 25
        34077 => X"14",  -- 20
        34078 => X"2A",  -- 42
        34079 => X"63",  -- 99
        34080 => X"8A",  -- 138
        34081 => X"AE",  -- 174
        34082 => X"BE",  -- 190
        34083 => X"B8",  -- 184
        34084 => X"B9",  -- 185
        34085 => X"C2",  -- 194
        34086 => X"C1",  -- 193
        34087 => X"BB",  -- 187
        34088 => X"CB",  -- 203
        34089 => X"C8",  -- 200
        34090 => X"C4",  -- 196
        34091 => X"BE",  -- 190
        34092 => X"BF",  -- 191
        34093 => X"BD",  -- 189
        34094 => X"AF",  -- 175
        34095 => X"9D",  -- 157
        34096 => X"A6",  -- 166
        34097 => X"95",  -- 149
        34098 => X"8F",  -- 143
        34099 => X"8C",  -- 140
        34100 => X"79",  -- 121
        34101 => X"5F",  -- 95
        34102 => X"4F",  -- 79
        34103 => X"43",  -- 67
        34104 => X"48",  -- 72
        34105 => X"2C",  -- 44
        34106 => X"18",  -- 24
        34107 => X"20",  -- 32
        34108 => X"3C",  -- 60
        34109 => X"5E",  -- 94
        34110 => X"71",  -- 113
        34111 => X"6F",  -- 111
        34112 => X"6A",  -- 106
        34113 => X"5E",  -- 94
        34114 => X"49",  -- 73
        34115 => X"33",  -- 51
        34116 => X"2C",  -- 44
        34117 => X"2C",  -- 44
        34118 => X"26",  -- 38
        34119 => X"1D",  -- 29
        34120 => X"2D",  -- 45
        34121 => X"44",  -- 68
        34122 => X"5C",  -- 92
        34123 => X"75",  -- 117
        34124 => X"92",  -- 146
        34125 => X"A2",  -- 162
        34126 => X"A4",  -- 164
        34127 => X"A5",  -- 165
        34128 => X"AE",  -- 174
        34129 => X"A8",  -- 168
        34130 => X"A1",  -- 161
        34131 => X"A3",  -- 163
        34132 => X"AD",  -- 173
        34133 => X"B3",  -- 179
        34134 => X"AC",  -- 172
        34135 => X"A2",  -- 162
        34136 => X"AA",  -- 170
        34137 => X"B0",  -- 176
        34138 => X"B5",  -- 181
        34139 => X"B5",  -- 181
        34140 => X"B9",  -- 185
        34141 => X"BD",  -- 189
        34142 => X"B8",  -- 184
        34143 => X"AE",  -- 174
        34144 => X"A2",  -- 162
        34145 => X"A5",  -- 165
        34146 => X"A7",  -- 167
        34147 => X"A8",  -- 168
        34148 => X"A7",  -- 167
        34149 => X"AA",  -- 170
        34150 => X"AD",  -- 173
        34151 => X"AF",  -- 175
        34152 => X"AC",  -- 172
        34153 => X"AE",  -- 174
        34154 => X"AD",  -- 173
        34155 => X"A9",  -- 169
        34156 => X"A6",  -- 166
        34157 => X"A2",  -- 162
        34158 => X"99",  -- 153
        34159 => X"90",  -- 144
        34160 => X"7F",  -- 127
        34161 => X"72",  -- 114
        34162 => X"59",  -- 89
        34163 => X"39",  -- 57
        34164 => X"26",  -- 38
        34165 => X"2A",  -- 42
        34166 => X"41",  -- 65
        34167 => X"55",  -- 85
        34168 => X"56",  -- 86
        34169 => X"6D",  -- 109
        34170 => X"69",  -- 105
        34171 => X"5F",  -- 95
        34172 => X"5D",  -- 93
        34173 => X"6D",  -- 109
        34174 => X"83",  -- 131
        34175 => X"7F",  -- 127
        34176 => X"8B",  -- 139
        34177 => X"9A",  -- 154
        34178 => X"94",  -- 148
        34179 => X"8A",  -- 138
        34180 => X"90",  -- 144
        34181 => X"8C",  -- 140
        34182 => X"81",  -- 129
        34183 => X"84",  -- 132
        34184 => X"9E",  -- 158
        34185 => X"95",  -- 149
        34186 => X"96",  -- 150
        34187 => X"9A",  -- 154
        34188 => X"8F",  -- 143
        34189 => X"8C",  -- 140
        34190 => X"7A",  -- 122
        34191 => X"7C",  -- 124
        34192 => X"89",  -- 137
        34193 => X"92",  -- 146
        34194 => X"92",  -- 146
        34195 => X"80",  -- 128
        34196 => X"87",  -- 135
        34197 => X"70",  -- 112
        34198 => X"7C",  -- 124
        34199 => X"76",  -- 118
        34200 => X"7A",  -- 122
        34201 => X"75",  -- 117
        34202 => X"7B",  -- 123
        34203 => X"8A",  -- 138
        34204 => X"90",  -- 144
        34205 => X"8D",  -- 141
        34206 => X"93",  -- 147
        34207 => X"A0",  -- 160
        34208 => X"9B",  -- 155
        34209 => X"9F",  -- 159
        34210 => X"A2",  -- 162
        34211 => X"A3",  -- 163
        34212 => X"A8",  -- 168
        34213 => X"AE",  -- 174
        34214 => X"B3",  -- 179
        34215 => X"B5",  -- 181
        34216 => X"B2",  -- 178
        34217 => X"C0",  -- 192
        34218 => X"BA",  -- 186
        34219 => X"93",  -- 147
        34220 => X"77",  -- 119
        34221 => X"8A",  -- 138
        34222 => X"AA",  -- 170
        34223 => X"B8",  -- 184
        34224 => X"BD",  -- 189
        34225 => X"C0",  -- 192
        34226 => X"C4",  -- 196
        34227 => X"C8",  -- 200
        34228 => X"CE",  -- 206
        34229 => X"D3",  -- 211
        34230 => X"D0",  -- 208
        34231 => X"CB",  -- 203
        34232 => X"C0",  -- 192
        34233 => X"BD",  -- 189
        34234 => X"B8",  -- 184
        34235 => X"B8",  -- 184
        34236 => X"B6",  -- 182
        34237 => X"AD",  -- 173
        34238 => X"9F",  -- 159
        34239 => X"95",  -- 149
        34240 => X"51",  -- 81
        34241 => X"54",  -- 84
        34242 => X"57",  -- 87
        34243 => X"58",  -- 88
        34244 => X"59",  -- 89
        34245 => X"59",  -- 89
        34246 => X"5B",  -- 91
        34247 => X"5D",  -- 93
        34248 => X"62",  -- 98
        34249 => X"5F",  -- 95
        34250 => X"5E",  -- 94
        34251 => X"5F",  -- 95
        34252 => X"62",  -- 98
        34253 => X"61",  -- 97
        34254 => X"5E",  -- 94
        34255 => X"5A",  -- 90
        34256 => X"56",  -- 86
        34257 => X"50",  -- 80
        34258 => X"4C",  -- 76
        34259 => X"49",  -- 73
        34260 => X"4C",  -- 76
        34261 => X"4E",  -- 78
        34262 => X"52",  -- 82
        34263 => X"53",  -- 83
        34264 => X"4F",  -- 79
        34265 => X"4D",  -- 77
        34266 => X"52",  -- 82
        34267 => X"62",  -- 98
        34268 => X"6B",  -- 107
        34269 => X"6B",  -- 107
        34270 => X"6D",  -- 109
        34271 => X"70",  -- 112
        34272 => X"5C",  -- 92
        34273 => X"44",  -- 68
        34274 => X"26",  -- 38
        34275 => X"10",  -- 16
        34276 => X"10",  -- 16
        34277 => X"0C",  -- 12
        34278 => X"20",  -- 32
        34279 => X"62",  -- 98
        34280 => X"79",  -- 121
        34281 => X"7B",  -- 123
        34282 => X"53",  -- 83
        34283 => X"25",  -- 37
        34284 => X"12",  -- 18
        34285 => X"05",  -- 5
        34286 => X"1F",  -- 31
        34287 => X"5E",  -- 94
        34288 => X"84",  -- 132
        34289 => X"61",  -- 97
        34290 => X"24",  -- 36
        34291 => X"0D",  -- 13
        34292 => X"0F",  -- 15
        34293 => X"19",  -- 25
        34294 => X"46",  -- 70
        34295 => X"74",  -- 116
        34296 => X"99",  -- 153
        34297 => X"A2",  -- 162
        34298 => X"A9",  -- 169
        34299 => X"AA",  -- 170
        34300 => X"A7",  -- 167
        34301 => X"A2",  -- 162
        34302 => X"A0",  -- 160
        34303 => X"9D",  -- 157
        34304 => X"9E",  -- 158
        34305 => X"9D",  -- 157
        34306 => X"94",  -- 148
        34307 => X"90",  -- 144
        34308 => X"89",  -- 137
        34309 => X"6F",  -- 111
        34310 => X"56",  -- 86
        34311 => X"54",  -- 84
        34312 => X"62",  -- 98
        34313 => X"6E",  -- 110
        34314 => X"66",  -- 102
        34315 => X"59",  -- 89
        34316 => X"4E",  -- 78
        34317 => X"2B",  -- 43
        34318 => X"0C",  -- 12
        34319 => X"0E",  -- 14
        34320 => X"16",  -- 22
        34321 => X"5E",  -- 94
        34322 => X"7B",  -- 123
        34323 => X"5D",  -- 93
        34324 => X"50",  -- 80
        34325 => X"2F",  -- 47
        34326 => X"11",  -- 17
        34327 => X"2F",  -- 47
        34328 => X"1B",  -- 27
        34329 => X"31",  -- 49
        34330 => X"62",  -- 98
        34331 => X"5A",  -- 90
        34332 => X"60",  -- 96
        34333 => X"65",  -- 101
        34334 => X"59",  -- 89
        34335 => X"40",  -- 64
        34336 => X"54",  -- 84
        34337 => X"58",  -- 88
        34338 => X"48",  -- 72
        34339 => X"54",  -- 84
        34340 => X"24",  -- 36
        34341 => X"25",  -- 37
        34342 => X"62",  -- 98
        34343 => X"68",  -- 104
        34344 => X"52",  -- 82
        34345 => X"5D",  -- 93
        34346 => X"62",  -- 98
        34347 => X"63",  -- 99
        34348 => X"55",  -- 85
        34349 => X"13",  -- 19
        34350 => X"0F",  -- 15
        34351 => X"42",  -- 66
        34352 => X"50",  -- 80
        34353 => X"5D",  -- 93
        34354 => X"86",  -- 134
        34355 => X"8C",  -- 140
        34356 => X"85",  -- 133
        34357 => X"7C",  -- 124
        34358 => X"75",  -- 117
        34359 => X"9C",  -- 156
        34360 => X"9B",  -- 155
        34361 => X"93",  -- 147
        34362 => X"94",  -- 148
        34363 => X"87",  -- 135
        34364 => X"8D",  -- 141
        34365 => X"91",  -- 145
        34366 => X"81",  -- 129
        34367 => X"99",  -- 153
        34368 => X"90",  -- 144
        34369 => X"85",  -- 133
        34370 => X"A9",  -- 169
        34371 => X"D1",  -- 209
        34372 => X"C3",  -- 195
        34373 => X"C5",  -- 197
        34374 => X"BA",  -- 186
        34375 => X"70",  -- 112
        34376 => X"26",  -- 38
        34377 => X"31",  -- 49
        34378 => X"16",  -- 22
        34379 => X"14",  -- 20
        34380 => X"1D",  -- 29
        34381 => X"23",  -- 35
        34382 => X"6A",  -- 106
        34383 => X"BC",  -- 188
        34384 => X"AD",  -- 173
        34385 => X"63",  -- 99
        34386 => X"26",  -- 38
        34387 => X"1C",  -- 28
        34388 => X"1F",  -- 31
        34389 => X"43",  -- 67
        34390 => X"90",  -- 144
        34391 => X"BB",  -- 187
        34392 => X"8B",  -- 139
        34393 => X"50",  -- 80
        34394 => X"17",  -- 23
        34395 => X"0C",  -- 12
        34396 => X"15",  -- 21
        34397 => X"0C",  -- 12
        34398 => X"1C",  -- 28
        34399 => X"46",  -- 70
        34400 => X"85",  -- 133
        34401 => X"B0",  -- 176
        34402 => X"C4",  -- 196
        34403 => X"BB",  -- 187
        34404 => X"B9",  -- 185
        34405 => X"C2",  -- 194
        34406 => X"C8",  -- 200
        34407 => X"C9",  -- 201
        34408 => X"C8",  -- 200
        34409 => X"CD",  -- 205
        34410 => X"CC",  -- 204
        34411 => X"C2",  -- 194
        34412 => X"BB",  -- 187
        34413 => X"B5",  -- 181
        34414 => X"A8",  -- 168
        34415 => X"9C",  -- 156
        34416 => X"96",  -- 150
        34417 => X"93",  -- 147
        34418 => X"91",  -- 145
        34419 => X"86",  -- 134
        34420 => X"78",  -- 120
        34421 => X"6D",  -- 109
        34422 => X"56",  -- 86
        34423 => X"39",  -- 57
        34424 => X"27",  -- 39
        34425 => X"1E",  -- 30
        34426 => X"1D",  -- 29
        34427 => X"26",  -- 38
        34428 => X"3A",  -- 58
        34429 => X"5A",  -- 90
        34430 => X"6E",  -- 110
        34431 => X"6C",  -- 108
        34432 => X"5F",  -- 95
        34433 => X"60",  -- 96
        34434 => X"53",  -- 83
        34435 => X"37",  -- 55
        34436 => X"23",  -- 35
        34437 => X"21",  -- 33
        34438 => X"25",  -- 37
        34439 => X"26",  -- 38
        34440 => X"31",  -- 49
        34441 => X"50",  -- 80
        34442 => X"60",  -- 96
        34443 => X"6F",  -- 111
        34444 => X"92",  -- 146
        34445 => X"A6",  -- 166
        34446 => X"A6",  -- 166
        34447 => X"A4",  -- 164
        34448 => X"A3",  -- 163
        34449 => X"AA",  -- 170
        34450 => X"AA",  -- 170
        34451 => X"A3",  -- 163
        34452 => X"A1",  -- 161
        34453 => X"A5",  -- 165
        34454 => X"A7",  -- 167
        34455 => X"A6",  -- 166
        34456 => X"AF",  -- 175
        34457 => X"B1",  -- 177
        34458 => X"AF",  -- 175
        34459 => X"AA",  -- 170
        34460 => X"AA",  -- 170
        34461 => X"AE",  -- 174
        34462 => X"AF",  -- 175
        34463 => X"AC",  -- 172
        34464 => X"A2",  -- 162
        34465 => X"A4",  -- 164
        34466 => X"A7",  -- 167
        34467 => X"A8",  -- 168
        34468 => X"A6",  -- 166
        34469 => X"A3",  -- 163
        34470 => X"A4",  -- 164
        34471 => X"A4",  -- 164
        34472 => X"A4",  -- 164
        34473 => X"A6",  -- 166
        34474 => X"A9",  -- 169
        34475 => X"AA",  -- 170
        34476 => X"AB",  -- 171
        34477 => X"A5",  -- 165
        34478 => X"97",  -- 151
        34479 => X"8A",  -- 138
        34480 => X"7D",  -- 125
        34481 => X"6A",  -- 106
        34482 => X"4E",  -- 78
        34483 => X"33",  -- 51
        34484 => X"20",  -- 32
        34485 => X"23",  -- 35
        34486 => X"38",  -- 56
        34487 => X"4C",  -- 76
        34488 => X"55",  -- 85
        34489 => X"6D",  -- 109
        34490 => X"76",  -- 118
        34491 => X"79",  -- 121
        34492 => X"7B",  -- 123
        34493 => X"86",  -- 134
        34494 => X"9C",  -- 156
        34495 => X"9C",  -- 156
        34496 => X"A2",  -- 162
        34497 => X"A3",  -- 163
        34498 => X"97",  -- 151
        34499 => X"94",  -- 148
        34500 => X"9E",  -- 158
        34501 => X"9D",  -- 157
        34502 => X"8F",  -- 143
        34503 => X"86",  -- 134
        34504 => X"9D",  -- 157
        34505 => X"9C",  -- 156
        34506 => X"96",  -- 150
        34507 => X"98",  -- 152
        34508 => X"9C",  -- 156
        34509 => X"91",  -- 145
        34510 => X"7B",  -- 123
        34511 => X"80",  -- 128
        34512 => X"8A",  -- 138
        34513 => X"8E",  -- 142
        34514 => X"90",  -- 144
        34515 => X"71",  -- 113
        34516 => X"7B",  -- 123
        34517 => X"68",  -- 104
        34518 => X"7A",  -- 122
        34519 => X"78",  -- 120
        34520 => X"86",  -- 134
        34521 => X"7F",  -- 127
        34522 => X"81",  -- 129
        34523 => X"8E",  -- 142
        34524 => X"95",  -- 149
        34525 => X"92",  -- 146
        34526 => X"93",  -- 147
        34527 => X"9A",  -- 154
        34528 => X"97",  -- 151
        34529 => X"9B",  -- 155
        34530 => X"A1",  -- 161
        34531 => X"A7",  -- 167
        34532 => X"AD",  -- 173
        34533 => X"B4",  -- 180
        34534 => X"B4",  -- 180
        34535 => X"B1",  -- 177
        34536 => X"B5",  -- 181
        34537 => X"B8",  -- 184
        34538 => X"BD",  -- 189
        34539 => X"A6",  -- 166
        34540 => X"7B",  -- 123
        34541 => X"79",  -- 121
        34542 => X"9F",  -- 159
        34543 => X"B8",  -- 184
        34544 => X"C1",  -- 193
        34545 => X"C3",  -- 195
        34546 => X"C3",  -- 195
        34547 => X"C3",  -- 195
        34548 => X"C9",  -- 201
        34549 => X"CF",  -- 207
        34550 => X"CF",  -- 207
        34551 => X"CC",  -- 204
        34552 => X"C3",  -- 195
        34553 => X"BC",  -- 188
        34554 => X"B6",  -- 182
        34555 => X"B3",  -- 179
        34556 => X"B1",  -- 177
        34557 => X"A7",  -- 167
        34558 => X"9B",  -- 155
        34559 => X"93",  -- 147
        34560 => X"52",  -- 82
        34561 => X"54",  -- 84
        34562 => X"56",  -- 86
        34563 => X"55",  -- 85
        34564 => X"54",  -- 84
        34565 => X"53",  -- 83
        34566 => X"55",  -- 85
        34567 => X"57",  -- 87
        34568 => X"60",  -- 96
        34569 => X"60",  -- 96
        34570 => X"5F",  -- 95
        34571 => X"5F",  -- 95
        34572 => X"5D",  -- 93
        34573 => X"58",  -- 88
        34574 => X"53",  -- 83
        34575 => X"4E",  -- 78
        34576 => X"47",  -- 71
        34577 => X"45",  -- 69
        34578 => X"43",  -- 67
        34579 => X"44",  -- 68
        34580 => X"46",  -- 70
        34581 => X"4A",  -- 74
        34582 => X"4D",  -- 77
        34583 => X"4F",  -- 79
        34584 => X"51",  -- 81
        34585 => X"51",  -- 81
        34586 => X"5C",  -- 92
        34587 => X"6C",  -- 108
        34588 => X"72",  -- 114
        34589 => X"6F",  -- 111
        34590 => X"70",  -- 112
        34591 => X"74",  -- 116
        34592 => X"64",  -- 100
        34593 => X"4F",  -- 79
        34594 => X"2E",  -- 46
        34595 => X"0E",  -- 14
        34596 => X"0B",  -- 11
        34597 => X"0A",  -- 10
        34598 => X"20",  -- 32
        34599 => X"5E",  -- 94
        34600 => X"74",  -- 116
        34601 => X"77",  -- 119
        34602 => X"4E",  -- 78
        34603 => X"21",  -- 33
        34604 => X"0D",  -- 13
        34605 => X"04",  -- 4
        34606 => X"27",  -- 39
        34607 => X"73",  -- 115
        34608 => X"83",  -- 131
        34609 => X"6D",  -- 109
        34610 => X"39",  -- 57
        34611 => X"27",  -- 39
        34612 => X"2B",  -- 43
        34613 => X"25",  -- 37
        34614 => X"35",  -- 53
        34615 => X"4F",  -- 79
        34616 => X"6F",  -- 111
        34617 => X"61",  -- 97
        34618 => X"5E",  -- 94
        34619 => X"72",  -- 114
        34620 => X"89",  -- 137
        34621 => X"8A",  -- 138
        34622 => X"70",  -- 112
        34623 => X"54",  -- 84
        34624 => X"57",  -- 87
        34625 => X"4B",  -- 75
        34626 => X"3D",  -- 61
        34627 => X"45",  -- 69
        34628 => X"5F",  -- 95
        34629 => X"6E",  -- 110
        34630 => X"69",  -- 105
        34631 => X"61",  -- 97
        34632 => X"57",  -- 87
        34633 => X"60",  -- 96
        34634 => X"58",  -- 88
        34635 => X"4B",  -- 75
        34636 => X"45",  -- 69
        34637 => X"31",  -- 49
        34638 => X"13",  -- 19
        34639 => X"09",  -- 9
        34640 => X"26",  -- 38
        34641 => X"55",  -- 85
        34642 => X"60",  -- 96
        34643 => X"55",  -- 85
        34644 => X"40",  -- 64
        34645 => X"29",  -- 41
        34646 => X"2F",  -- 47
        34647 => X"39",  -- 57
        34648 => X"1D",  -- 29
        34649 => X"3B",  -- 59
        34650 => X"67",  -- 103
        34651 => X"57",  -- 87
        34652 => X"56",  -- 86
        34653 => X"59",  -- 89
        34654 => X"5B",  -- 91
        34655 => X"43",  -- 67
        34656 => X"55",  -- 85
        34657 => X"40",  -- 64
        34658 => X"29",  -- 41
        34659 => X"4E",  -- 78
        34660 => X"43",  -- 67
        34661 => X"20",  -- 32
        34662 => X"69",  -- 105
        34663 => X"70",  -- 112
        34664 => X"56",  -- 86
        34665 => X"59",  -- 89
        34666 => X"5D",  -- 93
        34667 => X"51",  -- 81
        34668 => X"4B",  -- 75
        34669 => X"10",  -- 16
        34670 => X"0E",  -- 14
        34671 => X"43",  -- 67
        34672 => X"52",  -- 82
        34673 => X"49",  -- 73
        34674 => X"70",  -- 112
        34675 => X"83",  -- 131
        34676 => X"7D",  -- 125
        34677 => X"7C",  -- 124
        34678 => X"62",  -- 98
        34679 => X"4A",  -- 74
        34680 => X"22",  -- 34
        34681 => X"1A",  -- 26
        34682 => X"1E",  -- 30
        34683 => X"1E",  -- 30
        34684 => X"36",  -- 54
        34685 => X"44",  -- 68
        34686 => X"39",  -- 57
        34687 => X"50",  -- 80
        34688 => X"6D",  -- 109
        34689 => X"4E",  -- 78
        34690 => X"58",  -- 88
        34691 => X"99",  -- 153
        34692 => X"B7",  -- 183
        34693 => X"A6",  -- 166
        34694 => X"85",  -- 133
        34695 => X"54",  -- 84
        34696 => X"42",  -- 66
        34697 => X"65",  -- 101
        34698 => X"47",  -- 71
        34699 => X"2A",  -- 42
        34700 => X"1D",  -- 29
        34701 => X"1C",  -- 28
        34702 => X"63",  -- 99
        34703 => X"B3",  -- 179
        34704 => X"AF",  -- 175
        34705 => X"65",  -- 101
        34706 => X"28",  -- 40
        34707 => X"24",  -- 36
        34708 => X"23",  -- 35
        34709 => X"44",  -- 68
        34710 => X"8C",  -- 140
        34711 => X"AB",  -- 171
        34712 => X"9B",  -- 155
        34713 => X"4A",  -- 74
        34714 => X"16",  -- 22
        34715 => X"14",  -- 20
        34716 => X"12",  -- 18
        34717 => X"0F",  -- 15
        34718 => X"21",  -- 33
        34719 => X"35",  -- 53
        34720 => X"6C",  -- 108
        34721 => X"9E",  -- 158
        34722 => X"BE",  -- 190
        34723 => X"BB",  -- 187
        34724 => X"B5",  -- 181
        34725 => X"BB",  -- 187
        34726 => X"C8",  -- 200
        34727 => X"D5",  -- 213
        34728 => X"CE",  -- 206
        34729 => X"D1",  -- 209
        34730 => X"CF",  -- 207
        34731 => X"C4",  -- 196
        34732 => X"BD",  -- 189
        34733 => X"B6",  -- 182
        34734 => X"AC",  -- 172
        34735 => X"9F",  -- 159
        34736 => X"88",  -- 136
        34737 => X"87",  -- 135
        34738 => X"84",  -- 132
        34739 => X"7D",  -- 125
        34740 => X"74",  -- 116
        34741 => X"71",  -- 113
        34742 => X"61",  -- 97
        34743 => X"46",  -- 70
        34744 => X"1A",  -- 26
        34745 => X"18",  -- 24
        34746 => X"20",  -- 32
        34747 => X"2B",  -- 43
        34748 => X"3E",  -- 62
        34749 => X"59",  -- 89
        34750 => X"65",  -- 101
        34751 => X"5C",  -- 92
        34752 => X"51",  -- 81
        34753 => X"55",  -- 85
        34754 => X"4F",  -- 79
        34755 => X"38",  -- 56
        34756 => X"22",  -- 34
        34757 => X"1D",  -- 29
        34758 => X"20",  -- 32
        34759 => X"23",  -- 35
        34760 => X"3F",  -- 63
        34761 => X"5F",  -- 95
        34762 => X"6D",  -- 109
        34763 => X"74",  -- 116
        34764 => X"90",  -- 144
        34765 => X"A3",  -- 163
        34766 => X"A3",  -- 163
        34767 => X"9F",  -- 159
        34768 => X"9F",  -- 159
        34769 => X"AB",  -- 171
        34770 => X"B0",  -- 176
        34771 => X"A7",  -- 167
        34772 => X"A1",  -- 161
        34773 => X"A5",  -- 165
        34774 => X"AC",  -- 172
        34775 => X"B0",  -- 176
        34776 => X"A1",  -- 161
        34777 => X"AC",  -- 172
        34778 => X"B5",  -- 181
        34779 => X"B1",  -- 177
        34780 => X"A7",  -- 167
        34781 => X"A0",  -- 160
        34782 => X"9E",  -- 158
        34783 => X"9E",  -- 158
        34784 => X"9C",  -- 156
        34785 => X"A1",  -- 161
        34786 => X"A6",  -- 166
        34787 => X"A6",  -- 166
        34788 => X"A1",  -- 161
        34789 => X"99",  -- 153
        34790 => X"95",  -- 149
        34791 => X"93",  -- 147
        34792 => X"90",  -- 144
        34793 => X"92",  -- 146
        34794 => X"96",  -- 150
        34795 => X"9C",  -- 156
        34796 => X"A3",  -- 163
        34797 => X"A7",  -- 167
        34798 => X"9F",  -- 159
        34799 => X"95",  -- 149
        34800 => X"8E",  -- 142
        34801 => X"71",  -- 113
        34802 => X"53",  -- 83
        34803 => X"41",  -- 65
        34804 => X"3A",  -- 58
        34805 => X"38",  -- 56
        34806 => X"4A",  -- 74
        34807 => X"5E",  -- 94
        34808 => X"6F",  -- 111
        34809 => X"80",  -- 128
        34810 => X"8B",  -- 139
        34811 => X"9B",  -- 155
        34812 => X"99",  -- 153
        34813 => X"93",  -- 147
        34814 => X"A3",  -- 163
        34815 => X"AC",  -- 172
        34816 => X"B2",  -- 178
        34817 => X"AA",  -- 170
        34818 => X"A4",  -- 164
        34819 => X"A6",  -- 166
        34820 => X"AD",  -- 173
        34821 => X"A7",  -- 167
        34822 => X"9C",  -- 156
        34823 => X"98",  -- 152
        34824 => X"9E",  -- 158
        34825 => X"A3",  -- 163
        34826 => X"99",  -- 153
        34827 => X"9A",  -- 154
        34828 => X"A6",  -- 166
        34829 => X"91",  -- 145
        34830 => X"82",  -- 130
        34831 => X"85",  -- 133
        34832 => X"87",  -- 135
        34833 => X"86",  -- 134
        34834 => X"8C",  -- 140
        34835 => X"69",  -- 105
        34836 => X"7B",  -- 123
        34837 => X"71",  -- 113
        34838 => X"81",  -- 129
        34839 => X"83",  -- 131
        34840 => X"85",  -- 133
        34841 => X"85",  -- 133
        34842 => X"86",  -- 134
        34843 => X"8C",  -- 140
        34844 => X"97",  -- 151
        34845 => X"9F",  -- 159
        34846 => X"9E",  -- 158
        34847 => X"97",  -- 151
        34848 => X"97",  -- 151
        34849 => X"99",  -- 153
        34850 => X"9C",  -- 156
        34851 => X"A2",  -- 162
        34852 => X"AC",  -- 172
        34853 => X"B4",  -- 180
        34854 => X"B3",  -- 179
        34855 => X"AC",  -- 172
        34856 => X"B0",  -- 176
        34857 => X"A7",  -- 167
        34858 => X"B6",  -- 182
        34859 => X"BC",  -- 188
        34860 => X"90",  -- 144
        34861 => X"73",  -- 115
        34862 => X"8D",  -- 141
        34863 => X"B4",  -- 180
        34864 => X"C8",  -- 200
        34865 => X"C8",  -- 200
        34866 => X"C5",  -- 197
        34867 => X"C4",  -- 196
        34868 => X"C7",  -- 199
        34869 => X"CD",  -- 205
        34870 => X"CD",  -- 205
        34871 => X"C9",  -- 201
        34872 => X"CA",  -- 202
        34873 => X"C0",  -- 192
        34874 => X"B6",  -- 182
        34875 => X"B0",  -- 176
        34876 => X"A7",  -- 167
        34877 => X"9A",  -- 154
        34878 => X"8F",  -- 143
        34879 => X"8B",  -- 139
        34880 => X"58",  -- 88
        34881 => X"58",  -- 88
        34882 => X"57",  -- 87
        34883 => X"52",  -- 82
        34884 => X"4F",  -- 79
        34885 => X"4D",  -- 77
        34886 => X"4E",  -- 78
        34887 => X"51",  -- 81
        34888 => X"52",  -- 82
        34889 => X"53",  -- 83
        34890 => X"54",  -- 84
        34891 => X"53",  -- 83
        34892 => X"51",  -- 81
        34893 => X"4C",  -- 76
        34894 => X"49",  -- 73
        34895 => X"46",  -- 70
        34896 => X"40",  -- 64
        34897 => X"40",  -- 64
        34898 => X"40",  -- 64
        34899 => X"41",  -- 65
        34900 => X"42",  -- 66
        34901 => X"43",  -- 67
        34902 => X"43",  -- 67
        34903 => X"44",  -- 68
        34904 => X"4E",  -- 78
        34905 => X"53",  -- 83
        34906 => X"5C",  -- 92
        34907 => X"6A",  -- 106
        34908 => X"73",  -- 115
        34909 => X"74",  -- 116
        34910 => X"73",  -- 115
        34911 => X"74",  -- 116
        34912 => X"72",  -- 114
        34913 => X"5B",  -- 91
        34914 => X"36",  -- 54
        34915 => X"11",  -- 17
        34916 => X"0B",  -- 11
        34917 => X"08",  -- 8
        34918 => X"1B",  -- 27
        34919 => X"58",  -- 88
        34920 => X"87",  -- 135
        34921 => X"80",  -- 128
        34922 => X"4C",  -- 76
        34923 => X"19",  -- 25
        34924 => X"07",  -- 7
        34925 => X"04",  -- 4
        34926 => X"2C",  -- 44
        34927 => X"78",  -- 120
        34928 => X"80",  -- 128
        34929 => X"79",  -- 121
        34930 => X"57",  -- 87
        34931 => X"49",  -- 73
        34932 => X"41",  -- 65
        34933 => X"29",  -- 41
        34934 => X"22",  -- 34
        34935 => X"28",  -- 40
        34936 => X"2D",  -- 45
        34937 => X"2A",  -- 42
        34938 => X"37",  -- 55
        34939 => X"55",  -- 85
        34940 => X"6C",  -- 108
        34941 => X"62",  -- 98
        34942 => X"3D",  -- 61
        34943 => X"1C",  -- 28
        34944 => X"1A",  -- 26
        34945 => X"15",  -- 21
        34946 => X"14",  -- 20
        34947 => X"1A",  -- 26
        34948 => X"30",  -- 48
        34949 => X"4A",  -- 74
        34950 => X"5B",  -- 91
        34951 => X"60",  -- 96
        34952 => X"64",  -- 100
        34953 => X"6A",  -- 106
        34954 => X"5E",  -- 94
        34955 => X"45",  -- 69
        34956 => X"34",  -- 52
        34957 => X"23",  -- 35
        34958 => X"10",  -- 16
        34959 => X"07",  -- 7
        34960 => X"32",  -- 50
        34961 => X"46",  -- 70
        34962 => X"47",  -- 71
        34963 => X"4F",  -- 79
        34964 => X"3E",  -- 62
        34965 => X"34",  -- 52
        34966 => X"4D",  -- 77
        34967 => X"40",  -- 64
        34968 => X"3E",  -- 62
        34969 => X"56",  -- 86
        34970 => X"69",  -- 105
        34971 => X"55",  -- 85
        34972 => X"4C",  -- 76
        34973 => X"56",  -- 86
        34974 => X"5B",  -- 91
        34975 => X"46",  -- 70
        34976 => X"59",  -- 89
        34977 => X"41",  -- 65
        34978 => X"20",  -- 32
        34979 => X"24",  -- 36
        34980 => X"56",  -- 86
        34981 => X"42",  -- 66
        34982 => X"51",  -- 81
        34983 => X"6D",  -- 109
        34984 => X"55",  -- 85
        34985 => X"51",  -- 81
        34986 => X"5F",  -- 95
        34987 => X"4A",  -- 74
        34988 => X"46",  -- 70
        34989 => X"13",  -- 19
        34990 => X"13",  -- 19
        34991 => X"3F",  -- 63
        34992 => X"4B",  -- 75
        34993 => X"50",  -- 80
        34994 => X"7A",  -- 122
        34995 => X"9C",  -- 156
        34996 => X"83",  -- 131
        34997 => X"57",  -- 87
        34998 => X"32",  -- 50
        34999 => X"10",  -- 16
        35000 => X"1B",  -- 27
        35001 => X"1F",  -- 31
        35002 => X"23",  -- 35
        35003 => X"20",  -- 32
        35004 => X"30",  -- 48
        35005 => X"3B",  -- 59
        35006 => X"28",  -- 40
        35007 => X"1C",  -- 28
        35008 => X"1C",  -- 28
        35009 => X"47",  -- 71
        35010 => X"37",  -- 55
        35011 => X"3E",  -- 62
        35012 => X"7C",  -- 124
        35013 => X"81",  -- 129
        35014 => X"58",  -- 88
        35015 => X"41",  -- 65
        35016 => X"2C",  -- 44
        35017 => X"54",  -- 84
        35018 => X"72",  -- 114
        35019 => X"61",  -- 97
        35020 => X"2B",  -- 43
        35021 => X"21",  -- 33
        35022 => X"6F",  -- 111
        35023 => X"BC",  -- 188
        35024 => X"C3",  -- 195
        35025 => X"76",  -- 118
        35026 => X"2A",  -- 42
        35027 => X"25",  -- 37
        35028 => X"2A",  -- 42
        35029 => X"49",  -- 73
        35030 => X"8F",  -- 143
        35031 => X"A2",  -- 162
        35032 => X"B3",  -- 179
        35033 => X"52",  -- 82
        35034 => X"17",  -- 23
        35035 => X"17",  -- 23
        35036 => X"12",  -- 18
        35037 => X"16",  -- 22
        35038 => X"30",  -- 48
        35039 => X"41",  -- 65
        35040 => X"61",  -- 97
        35041 => X"92",  -- 146
        35042 => X"BA",  -- 186
        35043 => X"C2",  -- 194
        35044 => X"BD",  -- 189
        35045 => X"B7",  -- 183
        35046 => X"BD",  -- 189
        35047 => X"CB",  -- 203
        35048 => X"D5",  -- 213
        35049 => X"D1",  -- 209
        35050 => X"CA",  -- 202
        35051 => X"C4",  -- 196
        35052 => X"C3",  -- 195
        35053 => X"C1",  -- 193
        35054 => X"B3",  -- 179
        35055 => X"A1",  -- 161
        35056 => X"92",  -- 146
        35057 => X"7F",  -- 127
        35058 => X"78",  -- 120
        35059 => X"7A",  -- 122
        35060 => X"70",  -- 112
        35061 => X"62",  -- 98
        35062 => X"57",  -- 87
        35063 => X"4D",  -- 77
        35064 => X"2F",  -- 47
        35065 => X"24",  -- 36
        35066 => X"22",  -- 34
        35067 => X"2F",  -- 47
        35068 => X"46",  -- 70
        35069 => X"5B",  -- 91
        35070 => X"5A",  -- 90
        35071 => X"46",  -- 70
        35072 => X"41",  -- 65
        35073 => X"3C",  -- 60
        35074 => X"36",  -- 54
        35075 => X"2C",  -- 44
        35076 => X"22",  -- 34
        35077 => X"1D",  -- 29
        35078 => X"1B",  -- 27
        35079 => X"1B",  -- 27
        35080 => X"4A",  -- 74
        35081 => X"67",  -- 103
        35082 => X"7A",  -- 122
        35083 => X"7D",  -- 125
        35084 => X"89",  -- 137
        35085 => X"98",  -- 152
        35086 => X"98",  -- 152
        35087 => X"92",  -- 146
        35088 => X"9B",  -- 155
        35089 => X"A0",  -- 160
        35090 => X"A3",  -- 163
        35091 => X"A1",  -- 161
        35092 => X"A3",  -- 163
        35093 => X"A8",  -- 168
        35094 => X"AD",  -- 173
        35095 => X"B0",  -- 176
        35096 => X"AC",  -- 172
        35097 => X"A7",  -- 167
        35098 => X"A5",  -- 165
        35099 => X"A8",  -- 168
        35100 => X"AD",  -- 173
        35101 => X"AB",  -- 171
        35102 => X"9E",  -- 158
        35103 => X"91",  -- 145
        35104 => X"93",  -- 147
        35105 => X"99",  -- 153
        35106 => X"A0",  -- 160
        35107 => X"A2",  -- 162
        35108 => X"9E",  -- 158
        35109 => X"99",  -- 153
        35110 => X"95",  -- 149
        35111 => X"94",  -- 148
        35112 => X"8C",  -- 140
        35113 => X"8B",  -- 139
        35114 => X"88",  -- 136
        35115 => X"89",  -- 137
        35116 => X"91",  -- 145
        35117 => X"98",  -- 152
        35118 => X"97",  -- 151
        35119 => X"90",  -- 144
        35120 => X"84",  -- 132
        35121 => X"62",  -- 98
        35122 => X"47",  -- 71
        35123 => X"42",  -- 66
        35124 => X"47",  -- 71
        35125 => X"4F",  -- 79
        35126 => X"62",  -- 98
        35127 => X"77",  -- 119
        35128 => X"8C",  -- 140
        35129 => X"95",  -- 149
        35130 => X"9C",  -- 156
        35131 => X"AA",  -- 170
        35132 => X"A6",  -- 166
        35133 => X"96",  -- 150
        35134 => X"A3",  -- 163
        35135 => X"AF",  -- 175
        35136 => X"B1",  -- 177
        35137 => X"AF",  -- 175
        35138 => X"B2",  -- 178
        35139 => X"B6",  -- 182
        35140 => X"AF",  -- 175
        35141 => X"A5",  -- 165
        35142 => X"A4",  -- 164
        35143 => X"A9",  -- 169
        35144 => X"A3",  -- 163
        35145 => X"A6",  -- 166
        35146 => X"9B",  -- 155
        35147 => X"9B",  -- 155
        35148 => X"A5",  -- 165
        35149 => X"8B",  -- 139
        35150 => X"84",  -- 132
        35151 => X"83",  -- 131
        35152 => X"7D",  -- 125
        35153 => X"7D",  -- 125
        35154 => X"86",  -- 134
        35155 => X"6D",  -- 109
        35156 => X"83",  -- 131
        35157 => X"86",  -- 134
        35158 => X"8A",  -- 138
        35159 => X"8B",  -- 139
        35160 => X"8A",  -- 138
        35161 => X"91",  -- 145
        35162 => X"91",  -- 145
        35163 => X"8E",  -- 142
        35164 => X"97",  -- 151
        35165 => X"A4",  -- 164
        35166 => X"A0",  -- 160
        35167 => X"90",  -- 144
        35168 => X"9A",  -- 154
        35169 => X"9B",  -- 155
        35170 => X"9A",  -- 154
        35171 => X"9C",  -- 156
        35172 => X"A4",  -- 164
        35173 => X"B0",  -- 176
        35174 => X"B2",  -- 178
        35175 => X"B0",  -- 176
        35176 => X"A7",  -- 167
        35177 => X"97",  -- 151
        35178 => X"A6",  -- 166
        35179 => X"BD",  -- 189
        35180 => X"A5",  -- 165
        35181 => X"7E",  -- 126
        35182 => X"86",  -- 134
        35183 => X"AB",  -- 171
        35184 => X"CB",  -- 203
        35185 => X"CC",  -- 204
        35186 => X"CB",  -- 203
        35187 => X"C8",  -- 200
        35188 => X"C8",  -- 200
        35189 => X"CB",  -- 203
        35190 => X"CD",  -- 205
        35191 => X"CC",  -- 204
        35192 => X"CC",  -- 204
        35193 => X"C1",  -- 193
        35194 => X"B8",  -- 184
        35195 => X"AE",  -- 174
        35196 => X"A0",  -- 160
        35197 => X"8D",  -- 141
        35198 => X"81",  -- 129
        35199 => X"80",  -- 128
        35200 => X"5F",  -- 95
        35201 => X"5D",  -- 93
        35202 => X"5A",  -- 90
        35203 => X"54",  -- 84
        35204 => X"50",  -- 80
        35205 => X"4F",  -- 79
        35206 => X"52",  -- 82
        35207 => X"55",  -- 85
        35208 => X"53",  -- 83
        35209 => X"53",  -- 83
        35210 => X"52",  -- 82
        35211 => X"4E",  -- 78
        35212 => X"49",  -- 73
        35213 => X"46",  -- 70
        35214 => X"45",  -- 69
        35215 => X"45",  -- 69
        35216 => X"44",  -- 68
        35217 => X"45",  -- 69
        35218 => X"45",  -- 69
        35219 => X"44",  -- 68
        35220 => X"41",  -- 65
        35221 => X"3E",  -- 62
        35222 => X"3C",  -- 60
        35223 => X"3C",  -- 60
        35224 => X"43",  -- 67
        35225 => X"47",  -- 71
        35226 => X"50",  -- 80
        35227 => X"5E",  -- 94
        35228 => X"70",  -- 112
        35229 => X"7E",  -- 126
        35230 => X"7F",  -- 127
        35231 => X"7A",  -- 122
        35232 => X"79",  -- 121
        35233 => X"5B",  -- 91
        35234 => X"33",  -- 51
        35235 => X"18",  -- 24
        35236 => X"12",  -- 18
        35237 => X"0A",  -- 10
        35238 => X"1B",  -- 27
        35239 => X"5D",  -- 93
        35240 => X"97",  -- 151
        35241 => X"89",  -- 137
        35242 => X"4A",  -- 74
        35243 => X"14",  -- 20
        35244 => X"0A",  -- 10
        35245 => X"0B",  -- 11
        35246 => X"2F",  -- 47
        35247 => X"73",  -- 115
        35248 => X"81",  -- 129
        35249 => X"81",  -- 129
        35250 => X"6D",  -- 109
        35251 => X"5D",  -- 93
        35252 => X"48",  -- 72
        35253 => X"2C",  -- 44
        35254 => X"2A",  -- 42
        35255 => X"30",  -- 48
        35256 => X"2A",  -- 42
        35257 => X"2E",  -- 46
        35258 => X"3B",  -- 59
        35259 => X"44",  -- 68
        35260 => X"3E",  -- 62
        35261 => X"2C",  -- 44
        35262 => X"23",  -- 35
        35263 => X"23",  -- 35
        35264 => X"2B",  -- 43
        35265 => X"2C",  -- 44
        35266 => X"2A",  -- 42
        35267 => X"1D",  -- 29
        35268 => X"0F",  -- 15
        35269 => X"16",  -- 22
        35270 => X"27",  -- 39
        35271 => X"31",  -- 49
        35272 => X"5B",  -- 91
        35273 => X"70",  -- 112
        35274 => X"75",  -- 117
        35275 => X"58",  -- 88
        35276 => X"35",  -- 53
        35277 => X"1E",  -- 30
        35278 => X"15",  -- 21
        35279 => X"14",  -- 20
        35280 => X"2B",  -- 43
        35281 => X"31",  -- 49
        35282 => X"3A",  -- 58
        35283 => X"43",  -- 67
        35284 => X"42",  -- 66
        35285 => X"47",  -- 71
        35286 => X"51",  -- 81
        35287 => X"4D",  -- 77
        35288 => X"54",  -- 84
        35289 => X"63",  -- 99
        35290 => X"64",  -- 100
        35291 => X"5B",  -- 91
        35292 => X"49",  -- 73
        35293 => X"50",  -- 80
        35294 => X"54",  -- 84
        35295 => X"4A",  -- 74
        35296 => X"5B",  -- 91
        35297 => X"54",  -- 84
        35298 => X"31",  -- 49
        35299 => X"21",  -- 33
        35300 => X"52",  -- 82
        35301 => X"58",  -- 88
        35302 => X"43",  -- 67
        35303 => X"60",  -- 96
        35304 => X"53",  -- 83
        35305 => X"46",  -- 70
        35306 => X"57",  -- 87
        35307 => X"3F",  -- 63
        35308 => X"43",  -- 67
        35309 => X"1F",  -- 31
        35310 => X"22",  -- 34
        35311 => X"41",  -- 65
        35312 => X"45",  -- 69
        35313 => X"78",  -- 120
        35314 => X"93",  -- 147
        35315 => X"A1",  -- 161
        35316 => X"74",  -- 116
        35317 => X"2A",  -- 42
        35318 => X"20",  -- 32
        35319 => X"26",  -- 38
        35320 => X"30",  -- 48
        35321 => X"33",  -- 51
        35322 => X"35",  -- 53
        35323 => X"42",  -- 66
        35324 => X"51",  -- 81
        35325 => X"58",  -- 88
        35326 => X"50",  -- 80
        35327 => X"32",  -- 50
        35328 => X"05",  -- 5
        35329 => X"25",  -- 37
        35330 => X"1A",  -- 26
        35331 => X"34",  -- 52
        35332 => X"69",  -- 105
        35333 => X"61",  -- 97
        35334 => X"4C",  -- 76
        35335 => X"59",  -- 89
        35336 => X"4E",  -- 78
        35337 => X"64",  -- 100
        35338 => X"97",  -- 151
        35339 => X"9E",  -- 158
        35340 => X"62",  -- 98
        35341 => X"2E",  -- 46
        35342 => X"4E",  -- 78
        35343 => X"A1",  -- 161
        35344 => X"C4",  -- 196
        35345 => X"7F",  -- 127
        35346 => X"29",  -- 41
        35347 => X"1D",  -- 29
        35348 => X"2A",  -- 42
        35349 => X"56",  -- 86
        35350 => X"AB",  -- 171
        35351 => X"C8",  -- 200
        35352 => X"B3",  -- 179
        35353 => X"57",  -- 87
        35354 => X"0F",  -- 15
        35355 => X"08",  -- 8
        35356 => X"0E",  -- 14
        35357 => X"12",  -- 18
        35358 => X"2A",  -- 42
        35359 => X"4B",  -- 75
        35360 => X"6E",  -- 110
        35361 => X"93",  -- 147
        35362 => X"B7",  -- 183
        35363 => X"C9",  -- 201
        35364 => X"CB",  -- 203
        35365 => X"BD",  -- 189
        35366 => X"B7",  -- 183
        35367 => X"C0",  -- 192
        35368 => X"CE",  -- 206
        35369 => X"CF",  -- 207
        35370 => X"CA",  -- 202
        35371 => X"C3",  -- 195
        35372 => X"C2",  -- 194
        35373 => X"BD",  -- 189
        35374 => X"AF",  -- 175
        35375 => X"9E",  -- 158
        35376 => X"9B",  -- 155
        35377 => X"86",  -- 134
        35378 => X"7E",  -- 126
        35379 => X"80",  -- 128
        35380 => X"74",  -- 116
        35381 => X"62",  -- 98
        35382 => X"50",  -- 80
        35383 => X"41",  -- 65
        35384 => X"3F",  -- 63
        35385 => X"2F",  -- 47
        35386 => X"2C",  -- 44
        35387 => X"3B",  -- 59
        35388 => X"4E",  -- 78
        35389 => X"5B",  -- 91
        35390 => X"53",  -- 83
        35391 => X"3E",  -- 62
        35392 => X"2C",  -- 44
        35393 => X"24",  -- 36
        35394 => X"21",  -- 33
        35395 => X"22",  -- 34
        35396 => X"1E",  -- 30
        35397 => X"1A",  -- 26
        35398 => X"1B",  -- 27
        35399 => X"23",  -- 35
        35400 => X"4C",  -- 76
        35401 => X"67",  -- 103
        35402 => X"85",  -- 133
        35403 => X"8D",  -- 141
        35404 => X"8B",  -- 139
        35405 => X"93",  -- 147
        35406 => X"98",  -- 152
        35407 => X"90",  -- 144
        35408 => X"96",  -- 150
        35409 => X"96",  -- 150
        35410 => X"98",  -- 152
        35411 => X"9C",  -- 156
        35412 => X"A0",  -- 160
        35413 => X"A1",  -- 161
        35414 => X"A4",  -- 164
        35415 => X"AA",  -- 170
        35416 => X"BA",  -- 186
        35417 => X"A9",  -- 169
        35418 => X"9B",  -- 155
        35419 => X"9E",  -- 158
        35420 => X"AA",  -- 170
        35421 => X"AE",  -- 174
        35422 => X"A4",  -- 164
        35423 => X"97",  -- 151
        35424 => X"90",  -- 144
        35425 => X"93",  -- 147
        35426 => X"98",  -- 152
        35427 => X"97",  -- 151
        35428 => X"95",  -- 149
        35429 => X"94",  -- 148
        35430 => X"95",  -- 149
        35431 => X"95",  -- 149
        35432 => X"8A",  -- 138
        35433 => X"88",  -- 136
        35434 => X"82",  -- 130
        35435 => X"7E",  -- 126
        35436 => X"7E",  -- 126
        35437 => X"7E",  -- 126
        35438 => X"7C",  -- 124
        35439 => X"76",  -- 118
        35440 => X"6A",  -- 106
        35441 => X"55",  -- 85
        35442 => X"42",  -- 66
        35443 => X"41",  -- 65
        35444 => X"50",  -- 80
        35445 => X"63",  -- 99
        35446 => X"76",  -- 118
        35447 => X"83",  -- 131
        35448 => X"98",  -- 152
        35449 => X"A0",  -- 160
        35450 => X"A5",  -- 165
        35451 => X"AF",  -- 175
        35452 => X"AA",  -- 170
        35453 => X"A1",  -- 161
        35454 => X"AD",  -- 173
        35455 => X"B4",  -- 180
        35456 => X"AF",  -- 175
        35457 => X"B4",  -- 180
        35458 => X"BB",  -- 187
        35459 => X"B8",  -- 184
        35460 => X"AD",  -- 173
        35461 => X"AA",  -- 170
        35462 => X"AD",  -- 173
        35463 => X"AB",  -- 171
        35464 => X"A6",  -- 166
        35465 => X"A7",  -- 167
        35466 => X"A0",  -- 160
        35467 => X"9C",  -- 156
        35468 => X"A3",  -- 163
        35469 => X"85",  -- 133
        35470 => X"8A",  -- 138
        35471 => X"85",  -- 133
        35472 => X"7D",  -- 125
        35473 => X"7D",  -- 125
        35474 => X"82",  -- 130
        35475 => X"73",  -- 115
        35476 => X"87",  -- 135
        35477 => X"97",  -- 151
        35478 => X"8F",  -- 143
        35479 => X"8E",  -- 142
        35480 => X"90",  -- 144
        35481 => X"9B",  -- 155
        35482 => X"9D",  -- 157
        35483 => X"96",  -- 150
        35484 => X"97",  -- 151
        35485 => X"9F",  -- 159
        35486 => X"9C",  -- 156
        35487 => X"90",  -- 144
        35488 => X"99",  -- 153
        35489 => X"9F",  -- 159
        35490 => X"A0",  -- 160
        35491 => X"A1",  -- 161
        35492 => X"A3",  -- 163
        35493 => X"AB",  -- 171
        35494 => X"B1",  -- 177
        35495 => X"B4",  -- 180
        35496 => X"A4",  -- 164
        35497 => X"95",  -- 149
        35498 => X"93",  -- 147
        35499 => X"A4",  -- 164
        35500 => X"A9",  -- 169
        35501 => X"93",  -- 147
        35502 => X"8D",  -- 141
        35503 => X"9E",  -- 158
        35504 => X"C6",  -- 198
        35505 => X"CA",  -- 202
        35506 => X"CE",  -- 206
        35507 => X"CB",  -- 203
        35508 => X"C9",  -- 201
        35509 => X"CC",  -- 204
        35510 => X"CF",  -- 207
        35511 => X"CF",  -- 207
        35512 => X"CA",  -- 202
        35513 => X"C5",  -- 197
        35514 => X"BD",  -- 189
        35515 => X"B1",  -- 177
        35516 => X"9B",  -- 155
        35517 => X"81",  -- 129
        35518 => X"73",  -- 115
        35519 => X"73",  -- 115
        35520 => X"61",  -- 97
        35521 => X"60",  -- 96
        35522 => X"5D",  -- 93
        35523 => X"57",  -- 87
        35524 => X"55",  -- 85
        35525 => X"56",  -- 86
        35526 => X"5B",  -- 91
        35527 => X"5F",  -- 95
        35528 => X"65",  -- 101
        35529 => X"62",  -- 98
        35530 => X"5D",  -- 93
        35531 => X"55",  -- 85
        35532 => X"4E",  -- 78
        35533 => X"4A",  -- 74
        35534 => X"4A",  -- 74
        35535 => X"4A",  -- 74
        35536 => X"47",  -- 71
        35537 => X"49",  -- 73
        35538 => X"49",  -- 73
        35539 => X"47",  -- 71
        35540 => X"45",  -- 69
        35541 => X"40",  -- 64
        35542 => X"3C",  -- 60
        35543 => X"3B",  -- 59
        35544 => X"38",  -- 56
        35545 => X"3A",  -- 58
        35546 => X"41",  -- 65
        35547 => X"52",  -- 82
        35548 => X"6D",  -- 109
        35549 => X"87",  -- 135
        35550 => X"8A",  -- 138
        35551 => X"80",  -- 128
        35552 => X"78",  -- 120
        35553 => X"4F",  -- 79
        35554 => X"2A",  -- 42
        35555 => X"18",  -- 24
        35556 => X"17",  -- 23
        35557 => X"07",  -- 7
        35558 => X"1A",  -- 26
        35559 => X"64",  -- 100
        35560 => X"93",  -- 147
        35561 => X"82",  -- 130
        35562 => X"45",  -- 69
        35563 => X"14",  -- 20
        35564 => X"14",  -- 20
        35565 => X"1D",  -- 29
        35566 => X"3C",  -- 60
        35567 => X"73",  -- 115
        35568 => X"7D",  -- 125
        35569 => X"81",  -- 129
        35570 => X"72",  -- 114
        35571 => X"63",  -- 99
        35572 => X"4A",  -- 74
        35573 => X"3A",  -- 58
        35574 => X"4C",  -- 76
        35575 => X"5C",  -- 92
        35576 => X"6B",  -- 107
        35577 => X"56",  -- 86
        35578 => X"38",  -- 56
        35579 => X"1C",  -- 28
        35580 => X"09",  -- 9
        35581 => X"07",  -- 7
        35582 => X"22",  -- 34
        35583 => X"42",  -- 66
        35584 => X"3F",  -- 63
        35585 => X"33",  -- 51
        35586 => X"29",  -- 41
        35587 => X"1C",  -- 28
        35588 => X"0E",  -- 14
        35589 => X"10",  -- 16
        35590 => X"1A",  -- 26
        35591 => X"1B",  -- 27
        35592 => X"37",  -- 55
        35593 => X"64",  -- 100
        35594 => X"83",  -- 131
        35595 => X"73",  -- 115
        35596 => X"48",  -- 72
        35597 => X"2A",  -- 42
        35598 => X"27",  -- 39
        35599 => X"2B",  -- 43
        35600 => X"23",  -- 35
        35601 => X"25",  -- 37
        35602 => X"38",  -- 56
        35603 => X"38",  -- 56
        35604 => X"42",  -- 66
        35605 => X"52",  -- 82
        35606 => X"4A",  -- 74
        35607 => X"5B",  -- 91
        35608 => X"53",  -- 83
        35609 => X"61",  -- 97
        35610 => X"60",  -- 96
        35611 => X"68",  -- 104
        35612 => X"4C",  -- 76
        35613 => X"4C",  -- 76
        35614 => X"4F",  -- 79
        35615 => X"51",  -- 81
        35616 => X"56",  -- 86
        35617 => X"5D",  -- 93
        35618 => X"41",  -- 65
        35619 => X"44",  -- 68
        35620 => X"4A",  -- 74
        35621 => X"54",  -- 84
        35622 => X"4E",  -- 78
        35623 => X"5B",  -- 91
        35624 => X"55",  -- 85
        35625 => X"3E",  -- 62
        35626 => X"4D",  -- 77
        35627 => X"33",  -- 51
        35628 => X"3E",  -- 62
        35629 => X"27",  -- 39
        35630 => X"2F",  -- 47
        35631 => X"40",  -- 64
        35632 => X"4E",  -- 78
        35633 => X"A0",  -- 160
        35634 => X"97",  -- 151
        35635 => X"84",  -- 132
        35636 => X"5F",  -- 95
        35637 => X"1A",  -- 26
        35638 => X"29",  -- 41
        35639 => X"4D",  -- 77
        35640 => X"2C",  -- 44
        35641 => X"18",  -- 24
        35642 => X"0B",  -- 11
        35643 => X"2D",  -- 45
        35644 => X"41",  -- 65
        35645 => X"4A",  -- 74
        35646 => X"60",  -- 96
        35647 => X"53",  -- 83
        35648 => X"19",  -- 25
        35649 => X"00",  -- 0
        35650 => X"0A",  -- 10
        35651 => X"4F",  -- 79
        35652 => X"7A",  -- 122
        35653 => X"7C",  -- 124
        35654 => X"7C",  -- 124
        35655 => X"6F",  -- 111
        35656 => X"6F",  -- 111
        35657 => X"6B",  -- 107
        35658 => X"84",  -- 132
        35659 => X"A9",  -- 169
        35660 => X"B2",  -- 178
        35661 => X"6F",  -- 111
        35662 => X"57",  -- 87
        35663 => X"BD",  -- 189
        35664 => X"C4",  -- 196
        35665 => X"8D",  -- 141
        35666 => X"38",  -- 56
        35667 => X"1F",  -- 31
        35668 => X"23",  -- 35
        35669 => X"4C",  -- 76
        35670 => X"A8",  -- 168
        35671 => X"CC",  -- 204
        35672 => X"BD",  -- 189
        35673 => X"70",  -- 112
        35674 => X"1C",  -- 28
        35675 => X"0A",  -- 10
        35676 => X"1C",  -- 28
        35677 => X"16",  -- 22
        35678 => X"24",  -- 36
        35679 => X"55",  -- 85
        35680 => X"77",  -- 119
        35681 => X"8F",  -- 143
        35682 => X"AC",  -- 172
        35683 => X"C8",  -- 200
        35684 => X"D3",  -- 211
        35685 => X"C7",  -- 199
        35686 => X"BD",  -- 189
        35687 => X"C2",  -- 194
        35688 => X"C1",  -- 193
        35689 => X"CC",  -- 204
        35690 => X"CE",  -- 206
        35691 => X"C5",  -- 197
        35692 => X"B7",  -- 183
        35693 => X"AE",  -- 174
        35694 => X"A4",  -- 164
        35695 => X"9B",  -- 155
        35696 => X"91",  -- 145
        35697 => X"8C",  -- 140
        35698 => X"89",  -- 137
        35699 => X"85",  -- 133
        35700 => X"7D",  -- 125
        35701 => X"75",  -- 117
        35702 => X"5A",  -- 90
        35703 => X"35",  -- 53
        35704 => X"3B",  -- 59
        35705 => X"32",  -- 50
        35706 => X"37",  -- 55
        35707 => X"48",  -- 72
        35708 => X"53",  -- 83
        35709 => X"58",  -- 88
        35710 => X"51",  -- 81
        35711 => X"42",  -- 66
        35712 => X"1B",  -- 27
        35713 => X"19",  -- 25
        35714 => X"1C",  -- 28
        35715 => X"20",  -- 32
        35716 => X"19",  -- 25
        35717 => X"13",  -- 19
        35718 => X"1F",  -- 31
        35719 => X"35",  -- 53
        35720 => X"4D",  -- 77
        35721 => X"67",  -- 103
        35722 => X"8E",  -- 142
        35723 => X"9C",  -- 156
        35724 => X"95",  -- 149
        35725 => X"9B",  -- 155
        35726 => X"A5",  -- 165
        35727 => X"9C",  -- 156
        35728 => X"95",  -- 149
        35729 => X"96",  -- 150
        35730 => X"9D",  -- 157
        35731 => X"A0",  -- 160
        35732 => X"9B",  -- 155
        35733 => X"95",  -- 149
        35734 => X"9C",  -- 156
        35735 => X"A9",  -- 169
        35736 => X"AB",  -- 171
        35737 => X"AF",  -- 175
        35738 => X"B1",  -- 177
        35739 => X"AB",  -- 171
        35740 => X"A1",  -- 161
        35741 => X"9B",  -- 155
        35742 => X"A0",  -- 160
        35743 => X"A7",  -- 167
        35744 => X"95",  -- 149
        35745 => X"95",  -- 149
        35746 => X"91",  -- 145
        35747 => X"8A",  -- 138
        35748 => X"85",  -- 133
        35749 => X"84",  -- 132
        35750 => X"86",  -- 134
        35751 => X"89",  -- 137
        35752 => X"7C",  -- 124
        35753 => X"7D",  -- 125
        35754 => X"7A",  -- 122
        35755 => X"76",  -- 118
        35756 => X"71",  -- 113
        35757 => X"6E",  -- 110
        35758 => X"67",  -- 103
        35759 => X"5D",  -- 93
        35760 => X"64",  -- 100
        35761 => X"5E",  -- 94
        35762 => X"54",  -- 84
        35763 => X"51",  -- 81
        35764 => X"62",  -- 98
        35765 => X"7B",  -- 123
        35766 => X"8B",  -- 139
        35767 => X"8D",  -- 141
        35768 => X"99",  -- 153
        35769 => X"A9",  -- 169
        35770 => X"AE",  -- 174
        35771 => X"B4",  -- 180
        35772 => X"B1",  -- 177
        35773 => X"AB",  -- 171
        35774 => X"B5",  -- 181
        35775 => X"B4",  -- 180
        35776 => X"B6",  -- 182
        35777 => X"BB",  -- 187
        35778 => X"BD",  -- 189
        35779 => X"B5",  -- 181
        35780 => X"B0",  -- 176
        35781 => X"B8",  -- 184
        35782 => X"B6",  -- 182
        35783 => X"A6",  -- 166
        35784 => X"AA",  -- 170
        35785 => X"A8",  -- 168
        35786 => X"A2",  -- 162
        35787 => X"A0",  -- 160
        35788 => X"A3",  -- 163
        35789 => X"85",  -- 133
        35790 => X"92",  -- 146
        35791 => X"89",  -- 137
        35792 => X"87",  -- 135
        35793 => X"83",  -- 131
        35794 => X"81",  -- 129
        35795 => X"75",  -- 117
        35796 => X"86",  -- 134
        35797 => X"9E",  -- 158
        35798 => X"8F",  -- 143
        35799 => X"8E",  -- 142
        35800 => X"8D",  -- 141
        35801 => X"99",  -- 153
        35802 => X"A0",  -- 160
        35803 => X"9D",  -- 157
        35804 => X"9A",  -- 154
        35805 => X"9E",  -- 158
        35806 => X"9E",  -- 158
        35807 => X"9A",  -- 154
        35808 => X"94",  -- 148
        35809 => X"A1",  -- 161
        35810 => X"AA",  -- 170
        35811 => X"A9",  -- 169
        35812 => X"A6",  -- 166
        35813 => X"A8",  -- 168
        35814 => X"B0",  -- 176
        35815 => X"B5",  -- 181
        35816 => X"A5",  -- 165
        35817 => X"9C",  -- 156
        35818 => X"89",  -- 137
        35819 => X"8C",  -- 140
        35820 => X"A3",  -- 163
        35821 => X"A5",  -- 165
        35822 => X"96",  -- 150
        35823 => X"93",  -- 147
        35824 => X"BF",  -- 191
        35825 => X"C7",  -- 199
        35826 => X"CC",  -- 204
        35827 => X"CB",  -- 203
        35828 => X"C7",  -- 199
        35829 => X"CA",  -- 202
        35830 => X"CF",  -- 207
        35831 => X"D2",  -- 210
        35832 => X"D2",  -- 210
        35833 => X"CD",  -- 205
        35834 => X"C5",  -- 197
        35835 => X"B7",  -- 183
        35836 => X"99",  -- 153
        35837 => X"75",  -- 117
        35838 => X"61",  -- 97
        35839 => X"5F",  -- 95
        35840 => X"5A",  -- 90
        35841 => X"56",  -- 86
        35842 => X"50",  -- 80
        35843 => X"50",  -- 80
        35844 => X"56",  -- 86
        35845 => X"5A",  -- 90
        35846 => X"5E",  -- 94
        35847 => X"5D",  -- 93
        35848 => X"63",  -- 99
        35849 => X"64",  -- 100
        35850 => X"65",  -- 101
        35851 => X"60",  -- 96
        35852 => X"5A",  -- 90
        35853 => X"54",  -- 84
        35854 => X"53",  -- 83
        35855 => X"53",  -- 83
        35856 => X"51",  -- 81
        35857 => X"4F",  -- 79
        35858 => X"4C",  -- 76
        35859 => X"4C",  -- 76
        35860 => X"4A",  -- 74
        35861 => X"47",  -- 71
        35862 => X"41",  -- 65
        35863 => X"3D",  -- 61
        35864 => X"42",  -- 66
        35865 => X"2E",  -- 46
        35866 => X"3C",  -- 60
        35867 => X"67",  -- 103
        35868 => X"7F",  -- 127
        35869 => X"85",  -- 133
        35870 => X"8B",  -- 139
        35871 => X"94",  -- 148
        35872 => X"62",  -- 98
        35873 => X"52",  -- 82
        35874 => X"3C",  -- 60
        35875 => X"1F",  -- 31
        35876 => X"0E",  -- 14
        35877 => X"0D",  -- 13
        35878 => X"2C",  -- 44
        35879 => X"71",  -- 113
        35880 => X"84",  -- 132
        35881 => X"83",  -- 131
        35882 => X"4B",  -- 75
        35883 => X"11",  -- 17
        35884 => X"12",  -- 18
        35885 => X"09",  -- 9
        35886 => X"37",  -- 55
        35887 => X"75",  -- 117
        35888 => X"7E",  -- 126
        35889 => X"79",  -- 121
        35890 => X"6F",  -- 111
        35891 => X"4C",  -- 76
        35892 => X"44",  -- 68
        35893 => X"4B",  -- 75
        35894 => X"4D",  -- 77
        35895 => X"71",  -- 113
        35896 => X"92",  -- 146
        35897 => X"7C",  -- 124
        35898 => X"59",  -- 89
        35899 => X"29",  -- 41
        35900 => X"02",  -- 2
        35901 => X"02",  -- 2
        35902 => X"25",  -- 37
        35903 => X"4A",  -- 74
        35904 => X"47",  -- 71
        35905 => X"4B",  -- 75
        35906 => X"48",  -- 72
        35907 => X"3B",  -- 59
        35908 => X"2B",  -- 43
        35909 => X"28",  -- 40
        35910 => X"2E",  -- 46
        35911 => X"35",  -- 53
        35912 => X"1F",  -- 31
        35913 => X"41",  -- 65
        35914 => X"7F",  -- 127
        35915 => X"87",  -- 135
        35916 => X"67",  -- 103
        35917 => X"37",  -- 55
        35918 => X"2F",  -- 47
        35919 => X"21",  -- 33
        35920 => X"26",  -- 38
        35921 => X"2B",  -- 43
        35922 => X"2E",  -- 46
        35923 => X"33",  -- 51
        35924 => X"36",  -- 54
        35925 => X"32",  -- 50
        35926 => X"39",  -- 57
        35927 => X"4C",  -- 76
        35928 => X"4E",  -- 78
        35929 => X"54",  -- 84
        35930 => X"65",  -- 101
        35931 => X"61",  -- 97
        35932 => X"4A",  -- 74
        35933 => X"5D",  -- 93
        35934 => X"4B",  -- 75
        35935 => X"4F",  -- 79
        35936 => X"56",  -- 86
        35937 => X"4B",  -- 75
        35938 => X"49",  -- 73
        35939 => X"42",  -- 66
        35940 => X"54",  -- 84
        35941 => X"4C",  -- 76
        35942 => X"5A",  -- 90
        35943 => X"65",  -- 101
        35944 => X"55",  -- 85
        35945 => X"3B",  -- 59
        35946 => X"44",  -- 68
        35947 => X"3A",  -- 58
        35948 => X"3A",  -- 58
        35949 => X"2A",  -- 42
        35950 => X"37",  -- 55
        35951 => X"4A",  -- 74
        35952 => X"7F",  -- 127
        35953 => X"A9",  -- 169
        35954 => X"A8",  -- 168
        35955 => X"9C",  -- 156
        35956 => X"29",  -- 41
        35957 => X"1C",  -- 28
        35958 => X"79",  -- 121
        35959 => X"58",  -- 88
        35960 => X"53",  -- 83
        35961 => X"3B",  -- 59
        35962 => X"37",  -- 55
        35963 => X"55",  -- 85
        35964 => X"5B",  -- 91
        35965 => X"69",  -- 105
        35966 => X"7F",  -- 127
        35967 => X"61",  -- 97
        35968 => X"12",  -- 18
        35969 => X"14",  -- 20
        35970 => X"18",  -- 24
        35971 => X"64",  -- 100
        35972 => X"A9",  -- 169
        35973 => X"9A",  -- 154
        35974 => X"80",  -- 128
        35975 => X"6F",  -- 111
        35976 => X"59",  -- 89
        35977 => X"4E",  -- 78
        35978 => X"5C",  -- 92
        35979 => X"80",  -- 128
        35980 => X"B3",  -- 179
        35981 => X"A8",  -- 168
        35982 => X"7B",  -- 123
        35983 => X"92",  -- 146
        35984 => X"C4",  -- 196
        35985 => X"86",  -- 134
        35986 => X"38",  -- 56
        35987 => X"1F",  -- 31
        35988 => X"26",  -- 38
        35989 => X"6A",  -- 106
        35990 => X"B5",  -- 181
        35991 => X"D0",  -- 208
        35992 => X"BB",  -- 187
        35993 => X"71",  -- 113
        35994 => X"10",  -- 16
        35995 => X"16",  -- 22
        35996 => X"0C",  -- 12
        35997 => X"0F",  -- 15
        35998 => X"35",  -- 53
        35999 => X"4E",  -- 78
        36000 => X"6A",  -- 106
        36001 => X"92",  -- 146
        36002 => X"B5",  -- 181
        36003 => X"C2",  -- 194
        36004 => X"C9",  -- 201
        36005 => X"D0",  -- 208
        36006 => X"CA",  -- 202
        36007 => X"BB",  -- 187
        36008 => X"C3",  -- 195
        36009 => X"C6",  -- 198
        36010 => X"C6",  -- 198
        36011 => X"BE",  -- 190
        36012 => X"B0",  -- 176
        36013 => X"A5",  -- 165
        36014 => X"9E",  -- 158
        36015 => X"9D",  -- 157
        36016 => X"7B",  -- 123
        36017 => X"72",  -- 114
        36018 => X"71",  -- 113
        36019 => X"7C",  -- 124
        36020 => X"82",  -- 130
        36021 => X"77",  -- 119
        36022 => X"5E",  -- 94
        36023 => X"4A",  -- 74
        36024 => X"23",  -- 35
        36025 => X"33",  -- 51
        36026 => X"3B",  -- 59
        36027 => X"3C",  -- 60
        36028 => X"4E",  -- 78
        36029 => X"62",  -- 98
        36030 => X"52",  -- 82
        36031 => X"2E",  -- 46
        36032 => X"25",  -- 37
        36033 => X"1E",  -- 30
        36034 => X"17",  -- 23
        36035 => X"13",  -- 19
        36036 => X"15",  -- 21
        36037 => X"1E",  -- 30
        36038 => X"2C",  -- 44
        36039 => X"38",  -- 56
        36040 => X"5D",  -- 93
        36041 => X"7A",  -- 122
        36042 => X"8E",  -- 142
        36043 => X"95",  -- 149
        36044 => X"9B",  -- 155
        36045 => X"A0",  -- 160
        36046 => X"9E",  -- 158
        36047 => X"A0",  -- 160
        36048 => X"A4",  -- 164
        36049 => X"9E",  -- 158
        36050 => X"96",  -- 150
        36051 => X"99",  -- 153
        36052 => X"A1",  -- 161
        36053 => X"A4",  -- 164
        36054 => X"9B",  -- 155
        36055 => X"92",  -- 146
        36056 => X"9A",  -- 154
        36057 => X"A9",  -- 169
        36058 => X"B0",  -- 176
        36059 => X"AA",  -- 170
        36060 => X"9F",  -- 159
        36061 => X"9C",  -- 156
        36062 => X"99",  -- 153
        36063 => X"93",  -- 147
        36064 => X"A0",  -- 160
        36065 => X"98",  -- 152
        36066 => X"8B",  -- 139
        36067 => X"81",  -- 129
        36068 => X"7F",  -- 127
        36069 => X"81",  -- 129
        36070 => X"7A",  -- 122
        36071 => X"6E",  -- 110
        36072 => X"74",  -- 116
        36073 => X"73",  -- 115
        36074 => X"6F",  -- 111
        36075 => X"6A",  -- 106
        36076 => X"6A",  -- 106
        36077 => X"68",  -- 104
        36078 => X"5F",  -- 95
        36079 => X"52",  -- 82
        36080 => X"58",  -- 88
        36081 => X"62",  -- 98
        36082 => X"63",  -- 99
        36083 => X"71",  -- 113
        36084 => X"7A",  -- 122
        36085 => X"82",  -- 130
        36086 => X"98",  -- 152
        36087 => X"9F",  -- 159
        36088 => X"A8",  -- 168
        36089 => X"A3",  -- 163
        36090 => X"B9",  -- 185
        36091 => X"AE",  -- 174
        36092 => X"C0",  -- 192
        36093 => X"A8",  -- 168
        36094 => X"B8",  -- 184
        36095 => X"BA",  -- 186
        36096 => X"AE",  -- 174
        36097 => X"B4",  -- 180
        36098 => X"B0",  -- 176
        36099 => X"BB",  -- 187
        36100 => X"AF",  -- 175
        36101 => X"B5",  -- 181
        36102 => X"AF",  -- 175
        36103 => X"B6",  -- 182
        36104 => X"B7",  -- 183
        36105 => X"95",  -- 149
        36106 => X"9C",  -- 156
        36107 => X"A4",  -- 164
        36108 => X"92",  -- 146
        36109 => X"96",  -- 150
        36110 => X"78",  -- 120
        36111 => X"8D",  -- 141
        36112 => X"80",  -- 128
        36113 => X"81",  -- 129
        36114 => X"81",  -- 129
        36115 => X"7C",  -- 124
        36116 => X"79",  -- 121
        36117 => X"9D",  -- 157
        36118 => X"9C",  -- 156
        36119 => X"97",  -- 151
        36120 => X"96",  -- 150
        36121 => X"9F",  -- 159
        36122 => X"A1",  -- 161
        36123 => X"9B",  -- 155
        36124 => X"9C",  -- 156
        36125 => X"A4",  -- 164
        36126 => X"A8",  -- 168
        36127 => X"A6",  -- 166
        36128 => X"A1",  -- 161
        36129 => X"9E",  -- 158
        36130 => X"A7",  -- 167
        36131 => X"AA",  -- 170
        36132 => X"A7",  -- 167
        36133 => X"B3",  -- 179
        36134 => X"B6",  -- 182
        36135 => X"A4",  -- 164
        36136 => X"A6",  -- 166
        36137 => X"A1",  -- 161
        36138 => X"7E",  -- 126
        36139 => X"82",  -- 130
        36140 => X"92",  -- 146
        36141 => X"91",  -- 145
        36142 => X"9F",  -- 159
        36143 => X"A8",  -- 168
        36144 => X"AF",  -- 175
        36145 => X"C1",  -- 193
        36146 => X"CF",  -- 207
        36147 => X"CA",  -- 202
        36148 => X"C3",  -- 195
        36149 => X"C6",  -- 198
        36150 => X"CE",  -- 206
        36151 => X"D3",  -- 211
        36152 => X"CA",  -- 202
        36153 => X"D1",  -- 209
        36154 => X"C7",  -- 199
        36155 => X"B9",  -- 185
        36156 => X"A3",  -- 163
        36157 => X"79",  -- 121
        36158 => X"5B",  -- 91
        36159 => X"5D",  -- 93
        36160 => X"57",  -- 87
        36161 => X"53",  -- 83
        36162 => X"50",  -- 80
        36163 => X"51",  -- 81
        36164 => X"57",  -- 87
        36165 => X"5C",  -- 92
        36166 => X"5E",  -- 94
        36167 => X"5E",  -- 94
        36168 => X"5E",  -- 94
        36169 => X"5F",  -- 95
        36170 => X"5F",  -- 95
        36171 => X"5E",  -- 94
        36172 => X"5B",  -- 91
        36173 => X"59",  -- 89
        36174 => X"59",  -- 89
        36175 => X"59",  -- 89
        36176 => X"58",  -- 88
        36177 => X"55",  -- 85
        36178 => X"52",  -- 82
        36179 => X"50",  -- 80
        36180 => X"50",  -- 80
        36181 => X"4B",  -- 75
        36182 => X"45",  -- 69
        36183 => X"40",  -- 64
        36184 => X"3D",  -- 61
        36185 => X"39",  -- 57
        36186 => X"4E",  -- 78
        36187 => X"6F",  -- 111
        36188 => X"84",  -- 132
        36189 => X"89",  -- 137
        36190 => X"85",  -- 133
        36191 => X"7D",  -- 125
        36192 => X"65",  -- 101
        36193 => X"5C",  -- 92
        36194 => X"41",  -- 65
        36195 => X"18",  -- 24
        36196 => X"0B",  -- 11
        36197 => X"18",  -- 24
        36198 => X"34",  -- 52
        36199 => X"65",  -- 101
        36200 => X"8E",  -- 142
        36201 => X"86",  -- 134
        36202 => X"4C",  -- 76
        36203 => X"0E",  -- 14
        36204 => X"09",  -- 9
        36205 => X"07",  -- 7
        36206 => X"3F",  -- 63
        36207 => X"79",  -- 121
        36208 => X"6C",  -- 108
        36209 => X"66",  -- 102
        36210 => X"52",  -- 82
        36211 => X"2D",  -- 45
        36212 => X"28",  -- 40
        36213 => X"38",  -- 56
        36214 => X"49",  -- 73
        36215 => X"73",  -- 115
        36216 => X"A0",  -- 160
        36217 => X"B2",  -- 178
        36218 => X"79",  -- 121
        36219 => X"2C",  -- 44
        36220 => X"14",  -- 20
        36221 => X"09",  -- 9
        36222 => X"15",  -- 21
        36223 => X"46",  -- 70
        36224 => X"65",  -- 101
        36225 => X"5A",  -- 90
        36226 => X"4D",  -- 77
        36227 => X"47",  -- 71
        36228 => X"40",  -- 64
        36229 => X"3D",  -- 61
        36230 => X"47",  -- 71
        36231 => X"58",  -- 88
        36232 => X"13",  -- 19
        36233 => X"26",  -- 38
        36234 => X"66",  -- 102
        36235 => X"89",  -- 137
        36236 => X"7C",  -- 124
        36237 => X"45",  -- 69
        36238 => X"2D",  -- 45
        36239 => X"21",  -- 33
        36240 => X"28",  -- 40
        36241 => X"2C",  -- 44
        36242 => X"26",  -- 38
        36243 => X"22",  -- 34
        36244 => X"2A",  -- 42
        36245 => X"35",  -- 53
        36246 => X"3F",  -- 63
        36247 => X"4B",  -- 75
        36248 => X"51",  -- 81
        36249 => X"5A",  -- 90
        36250 => X"58",  -- 88
        36251 => X"61",  -- 97
        36252 => X"4F",  -- 79
        36253 => X"53",  -- 83
        36254 => X"51",  -- 81
        36255 => X"4B",  -- 75
        36256 => X"48",  -- 72
        36257 => X"43",  -- 67
        36258 => X"47",  -- 71
        36259 => X"47",  -- 71
        36260 => X"4D",  -- 77
        36261 => X"4E",  -- 78
        36262 => X"57",  -- 87
        36263 => X"5B",  -- 91
        36264 => X"52",  -- 82
        36265 => X"44",  -- 68
        36266 => X"50",  -- 80
        36267 => X"46",  -- 70
        36268 => X"40",  -- 64
        36269 => X"2D",  -- 45
        36270 => X"38",  -- 56
        36271 => X"55",  -- 85
        36272 => X"9C",  -- 156
        36273 => X"B6",  -- 182
        36274 => X"B2",  -- 178
        36275 => X"81",  -- 129
        36276 => X"1E",  -- 30
        36277 => X"1A",  -- 26
        36278 => X"74",  -- 116
        36279 => X"8F",  -- 143
        36280 => X"64",  -- 100
        36281 => X"60",  -- 96
        36282 => X"55",  -- 85
        36283 => X"5F",  -- 95
        36284 => X"74",  -- 116
        36285 => X"90",  -- 144
        36286 => X"88",  -- 136
        36287 => X"43",  -- 67
        36288 => X"09",  -- 9
        36289 => X"08",  -- 8
        36290 => X"49",  -- 73
        36291 => X"AD",  -- 173
        36292 => X"CE",  -- 206
        36293 => X"BA",  -- 186
        36294 => X"8F",  -- 143
        36295 => X"55",  -- 85
        36296 => X"2D",  -- 45
        36297 => X"2F",  -- 47
        36298 => X"47",  -- 71
        36299 => X"81",  -- 129
        36300 => X"C4",  -- 196
        36301 => X"C7",  -- 199
        36302 => X"97",  -- 151
        36303 => X"87",  -- 135
        36304 => X"B6",  -- 182
        36305 => X"8A",  -- 138
        36306 => X"43",  -- 67
        36307 => X"2B",  -- 43
        36308 => X"35",  -- 53
        36309 => X"80",  -- 128
        36310 => X"BE",  -- 190
        36311 => X"CA",  -- 202
        36312 => X"BE",  -- 190
        36313 => X"7A",  -- 122
        36314 => X"16",  -- 22
        36315 => X"11",  -- 17
        36316 => X"0A",  -- 10
        36317 => X"0D",  -- 13
        36318 => X"36",  -- 54
        36319 => X"5A",  -- 90
        36320 => X"79",  -- 121
        36321 => X"92",  -- 146
        36322 => X"AD",  -- 173
        36323 => X"BE",  -- 190
        36324 => X"C4",  -- 196
        36325 => X"C5",  -- 197
        36326 => X"C2",  -- 194
        36327 => X"BA",  -- 186
        36328 => X"C6",  -- 198
        36329 => X"CC",  -- 204
        36330 => X"CC",  -- 204
        36331 => X"C0",  -- 192
        36332 => X"AC",  -- 172
        36333 => X"98",  -- 152
        36334 => X"8C",  -- 140
        36335 => X"8A",  -- 138
        36336 => X"8C",  -- 140
        36337 => X"72",  -- 114
        36338 => X"5B",  -- 91
        36339 => X"5B",  -- 91
        36340 => X"67",  -- 103
        36341 => X"6A",  -- 106
        36342 => X"5F",  -- 95
        36343 => X"52",  -- 82
        36344 => X"3A",  -- 58
        36345 => X"22",  -- 34
        36346 => X"30",  -- 48
        36347 => X"40",  -- 64
        36348 => X"3C",  -- 60
        36349 => X"4C",  -- 76
        36350 => X"50",  -- 80
        36351 => X"2D",  -- 45
        36352 => X"1D",  -- 29
        36353 => X"1B",  -- 27
        36354 => X"1A",  -- 26
        36355 => X"1B",  -- 27
        36356 => X"1D",  -- 29
        36357 => X"27",  -- 39
        36358 => X"3C",  -- 60
        36359 => X"50",  -- 80
        36360 => X"67",  -- 103
        36361 => X"80",  -- 128
        36362 => X"91",  -- 145
        36363 => X"92",  -- 146
        36364 => X"97",  -- 151
        36365 => X"9A",  -- 154
        36366 => X"9C",  -- 156
        36367 => X"A2",  -- 162
        36368 => X"9F",  -- 159
        36369 => X"9E",  -- 158
        36370 => X"9E",  -- 158
        36371 => X"9E",  -- 158
        36372 => X"99",  -- 153
        36373 => X"94",  -- 148
        36374 => X"98",  -- 152
        36375 => X"A0",  -- 160
        36376 => X"A2",  -- 162
        36377 => X"A2",  -- 162
        36378 => X"A2",  -- 162
        36379 => X"A2",  -- 162
        36380 => X"9E",  -- 158
        36381 => X"98",  -- 152
        36382 => X"95",  -- 149
        36383 => X"94",  -- 148
        36384 => X"9C",  -- 156
        36385 => X"96",  -- 150
        36386 => X"89",  -- 137
        36387 => X"7A",  -- 122
        36388 => X"73",  -- 115
        36389 => X"71",  -- 113
        36390 => X"70",  -- 112
        36391 => X"6C",  -- 108
        36392 => X"6F",  -- 111
        36393 => X"6F",  -- 111
        36394 => X"6A",  -- 106
        36395 => X"63",  -- 99
        36396 => X"5E",  -- 94
        36397 => X"5B",  -- 91
        36398 => X"58",  -- 88
        36399 => X"52",  -- 82
        36400 => X"52",  -- 82
        36401 => X"66",  -- 102
        36402 => X"72",  -- 114
        36403 => X"83",  -- 131
        36404 => X"8B",  -- 139
        36405 => X"8E",  -- 142
        36406 => X"A1",  -- 161
        36407 => X"A6",  -- 166
        36408 => X"B2",  -- 178
        36409 => X"AC",  -- 172
        36410 => X"B7",  -- 183
        36411 => X"AE",  -- 174
        36412 => X"BC",  -- 188
        36413 => X"B2",  -- 178
        36414 => X"BE",  -- 190
        36415 => X"BF",  -- 191
        36416 => X"B3",  -- 179
        36417 => X"B8",  -- 184
        36418 => X"BC",  -- 188
        36419 => X"BF",  -- 191
        36420 => X"B4",  -- 180
        36421 => X"B3",  -- 179
        36422 => X"B3",  -- 179
        36423 => X"BD",  -- 189
        36424 => X"B5",  -- 181
        36425 => X"94",  -- 148
        36426 => X"A0",  -- 160
        36427 => X"A3",  -- 163
        36428 => X"96",  -- 150
        36429 => X"91",  -- 145
        36430 => X"7C",  -- 124
        36431 => X"8D",  -- 141
        36432 => X"85",  -- 133
        36433 => X"86",  -- 134
        36434 => X"88",  -- 136
        36435 => X"84",  -- 132
        36436 => X"7C",  -- 124
        36437 => X"9A",  -- 154
        36438 => X"97",  -- 151
        36439 => X"91",  -- 145
        36440 => X"A2",  -- 162
        36441 => X"97",  -- 151
        36442 => X"97",  -- 151
        36443 => X"A1",  -- 161
        36444 => X"A1",  -- 161
        36445 => X"97",  -- 151
        36446 => X"98",  -- 152
        36447 => X"A6",  -- 166
        36448 => X"A2",  -- 162
        36449 => X"A0",  -- 160
        36450 => X"A7",  -- 167
        36451 => X"A6",  -- 166
        36452 => X"A1",  -- 161
        36453 => X"AD",  -- 173
        36454 => X"B3",  -- 179
        36455 => X"A9",  -- 169
        36456 => X"A7",  -- 167
        36457 => X"A4",  -- 164
        36458 => X"84",  -- 132
        36459 => X"7A",  -- 122
        36460 => X"82",  -- 130
        36461 => X"8C",  -- 140
        36462 => X"AA",  -- 170
        36463 => X"B3",  -- 179
        36464 => X"B9",  -- 185
        36465 => X"BF",  -- 191
        36466 => X"C3",  -- 195
        36467 => X"C3",  -- 195
        36468 => X"C3",  -- 195
        36469 => X"C6",  -- 198
        36470 => X"C8",  -- 200
        36471 => X"C9",  -- 201
        36472 => X"D0",  -- 208
        36473 => X"D0",  -- 208
        36474 => X"C7",  -- 199
        36475 => X"BD",  -- 189
        36476 => X"A9",  -- 169
        36477 => X"7C",  -- 124
        36478 => X"5B",  -- 91
        36479 => X"5C",  -- 92
        36480 => X"57",  -- 87
        36481 => X"55",  -- 85
        36482 => X"53",  -- 83
        36483 => X"55",  -- 85
        36484 => X"5A",  -- 90
        36485 => X"5E",  -- 94
        36486 => X"5F",  -- 95
        36487 => X"5F",  -- 95
        36488 => X"5B",  -- 91
        36489 => X"5A",  -- 90
        36490 => X"59",  -- 89
        36491 => X"5A",  -- 90
        36492 => X"5B",  -- 91
        36493 => X"5C",  -- 92
        36494 => X"5C",  -- 92
        36495 => X"5B",  -- 91
        36496 => X"5C",  -- 92
        36497 => X"5A",  -- 90
        36498 => X"56",  -- 86
        36499 => X"56",  -- 86
        36500 => X"56",  -- 86
        36501 => X"52",  -- 82
        36502 => X"4C",  -- 76
        36503 => X"48",  -- 72
        36504 => X"41",  -- 65
        36505 => X"49",  -- 73
        36506 => X"5F",  -- 95
        36507 => X"75",  -- 117
        36508 => X"82",  -- 130
        36509 => X"8B",  -- 139
        36510 => X"83",  -- 131
        36511 => X"6D",  -- 109
        36512 => X"72",  -- 114
        36513 => X"63",  -- 99
        36514 => X"43",  -- 67
        36515 => X"19",  -- 25
        36516 => X"0F",  -- 15
        36517 => X"1D",  -- 29
        36518 => X"35",  -- 53
        36519 => X"62",  -- 98
        36520 => X"8E",  -- 142
        36521 => X"81",  -- 129
        36522 => X"4F",  -- 79
        36523 => X"13",  -- 19
        36524 => X"07",  -- 7
        36525 => X"0F",  -- 15
        36526 => X"53",  -- 83
        36527 => X"82",  -- 130
        36528 => X"82",  -- 130
        36529 => X"77",  -- 119
        36530 => X"54",  -- 84
        36531 => X"20",  -- 32
        36532 => X"11",  -- 17
        36533 => X"18",  -- 24
        36534 => X"28",  -- 40
        36535 => X"4D",  -- 77
        36536 => X"8D",  -- 141
        36537 => X"AD",  -- 173
        36538 => X"94",  -- 148
        36539 => X"48",  -- 72
        36540 => X"16",  -- 22
        36541 => X"08",  -- 8
        36542 => X"10",  -- 16
        36543 => X"23",  -- 35
        36544 => X"65",  -- 101
        36545 => X"71",  -- 113
        36546 => X"6B",  -- 107
        36547 => X"58",  -- 88
        36548 => X"56",  -- 86
        36549 => X"67",  -- 103
        36550 => X"69",  -- 105
        36551 => X"5C",  -- 92
        36552 => X"12",  -- 18
        36553 => X"0E",  -- 14
        36554 => X"43",  -- 67
        36555 => X"81",  -- 129
        36556 => X"96",  -- 150
        36557 => X"5C",  -- 92
        36558 => X"35",  -- 53
        36559 => X"28",  -- 40
        36560 => X"28",  -- 40
        36561 => X"2C",  -- 44
        36562 => X"22",  -- 34
        36563 => X"1B",  -- 27
        36564 => X"28",  -- 40
        36565 => X"3A",  -- 58
        36566 => X"43",  -- 67
        36567 => X"48",  -- 72
        36568 => X"57",  -- 87
        36569 => X"5B",  -- 91
        36570 => X"4C",  -- 76
        36571 => X"60",  -- 96
        36572 => X"54",  -- 84
        36573 => X"4C",  -- 76
        36574 => X"55",  -- 85
        36575 => X"48",  -- 72
        36576 => X"43",  -- 67
        36577 => X"42",  -- 66
        36578 => X"49",  -- 73
        36579 => X"52",  -- 82
        36580 => X"48",  -- 72
        36581 => X"53",  -- 83
        36582 => X"58",  -- 88
        36583 => X"50",  -- 80
        36584 => X"42",  -- 66
        36585 => X"45",  -- 69
        36586 => X"53",  -- 83
        36587 => X"47",  -- 71
        36588 => X"46",  -- 70
        36589 => X"36",  -- 54
        36590 => X"46",  -- 70
        36591 => X"74",  -- 116
        36592 => X"B2",  -- 178
        36593 => X"B3",  -- 179
        36594 => X"92",  -- 146
        36595 => X"3A",  -- 58
        36596 => X"04",  -- 4
        36597 => X"12",  -- 18
        36598 => X"58",  -- 88
        36599 => X"AC",  -- 172
        36600 => X"92",  -- 146
        36601 => X"8C",  -- 140
        36602 => X"7F",  -- 127
        36603 => X"8B",  -- 139
        36604 => X"A0",  -- 160
        36605 => X"99",  -- 153
        36606 => X"68",  -- 104
        36607 => X"23",  -- 35
        36608 => X"1F",  -- 31
        36609 => X"1D",  -- 29
        36610 => X"6F",  -- 111
        36611 => X"C5",  -- 197
        36612 => X"D4",  -- 212
        36613 => X"B6",  -- 182
        36614 => X"6F",  -- 111
        36615 => X"22",  -- 34
        36616 => X"0E",  -- 14
        36617 => X"12",  -- 18
        36618 => X"2B",  -- 43
        36619 => X"76",  -- 118
        36620 => X"B9",  -- 185
        36621 => X"CA",  -- 202
        36622 => X"C5",  -- 197
        36623 => X"BA",  -- 186
        36624 => X"B9",  -- 185
        36625 => X"92",  -- 146
        36626 => X"3F",  -- 63
        36627 => X"20",  -- 32
        36628 => X"2E",  -- 46
        36629 => X"89",  -- 137
        36630 => X"C9",  -- 201
        36631 => X"D1",  -- 209
        36632 => X"C9",  -- 201
        36633 => X"8E",  -- 142
        36634 => X"25",  -- 37
        36635 => X"0E",  -- 14
        36636 => X"0E",  -- 14
        36637 => X"12",  -- 18
        36638 => X"38",  -- 56
        36639 => X"68",  -- 104
        36640 => X"8B",  -- 139
        36641 => X"96",  -- 150
        36642 => X"A8",  -- 168
        36643 => X"B9",  -- 185
        36644 => X"BE",  -- 190
        36645 => X"BA",  -- 186
        36646 => X"B5",  -- 181
        36647 => X"B5",  -- 181
        36648 => X"C0",  -- 192
        36649 => X"CB",  -- 203
        36650 => X"D2",  -- 210
        36651 => X"C9",  -- 201
        36652 => X"B2",  -- 178
        36653 => X"9A",  -- 154
        36654 => X"8D",  -- 141
        36655 => X"88",  -- 136
        36656 => X"81",  -- 129
        36657 => X"72",  -- 114
        36658 => X"62",  -- 98
        36659 => X"55",  -- 85
        36660 => X"4D",  -- 77
        36661 => X"49",  -- 73
        36662 => X"4B",  -- 75
        36663 => X"4F",  -- 79
        36664 => X"48",  -- 72
        36665 => X"30",  -- 48
        36666 => X"3B",  -- 59
        36667 => X"48",  -- 72
        36668 => X"3B",  -- 59
        36669 => X"36",  -- 54
        36670 => X"3E",  -- 62
        36671 => X"3A",  -- 58
        36672 => X"1E",  -- 30
        36673 => X"1C",  -- 28
        36674 => X"20",  -- 32
        36675 => X"26",  -- 38
        36676 => X"29",  -- 41
        36677 => X"32",  -- 50
        36678 => X"4C",  -- 76
        36679 => X"68",  -- 104
        36680 => X"72",  -- 114
        36681 => X"87",  -- 135
        36682 => X"92",  -- 146
        36683 => X"8E",  -- 142
        36684 => X"8E",  -- 142
        36685 => X"91",  -- 145
        36686 => X"96",  -- 150
        36687 => X"A1",  -- 161
        36688 => X"A0",  -- 160
        36689 => X"9F",  -- 159
        36690 => X"9E",  -- 158
        36691 => X"9B",  -- 155
        36692 => X"92",  -- 146
        36693 => X"8B",  -- 139
        36694 => X"93",  -- 147
        36695 => X"A1",  -- 161
        36696 => X"A6",  -- 166
        36697 => X"9B",  -- 155
        36698 => X"98",  -- 152
        36699 => X"9E",  -- 158
        36700 => X"9F",  -- 159
        36701 => X"94",  -- 148
        36702 => X"8C",  -- 140
        36703 => X"8B",  -- 139
        36704 => X"89",  -- 137
        36705 => X"88",  -- 136
        36706 => X"82",  -- 130
        36707 => X"75",  -- 117
        36708 => X"69",  -- 105
        36709 => X"64",  -- 100
        36710 => X"63",  -- 99
        36711 => X"62",  -- 98
        36712 => X"5F",  -- 95
        36713 => X"61",  -- 97
        36714 => X"5C",  -- 92
        36715 => X"4F",  -- 79
        36716 => X"45",  -- 69
        36717 => X"44",  -- 68
        36718 => X"4B",  -- 75
        36719 => X"50",  -- 80
        36720 => X"56",  -- 86
        36721 => X"6F",  -- 111
        36722 => X"82",  -- 130
        36723 => X"95",  -- 149
        36724 => X"99",  -- 153
        36725 => X"98",  -- 152
        36726 => X"A8",  -- 168
        36727 => X"AD",  -- 173
        36728 => X"B7",  -- 183
        36729 => X"B7",  -- 183
        36730 => X"B5",  -- 181
        36731 => X"B4",  -- 180
        36732 => X"B9",  -- 185
        36733 => X"BE",  -- 190
        36734 => X"C1",  -- 193
        36735 => X"BE",  -- 190
        36736 => X"B3",  -- 179
        36737 => X"B6",  -- 182
        36738 => X"C1",  -- 193
        36739 => X"BC",  -- 188
        36740 => X"B5",  -- 181
        36741 => X"A9",  -- 169
        36742 => X"B0",  -- 176
        36743 => X"BA",  -- 186
        36744 => X"AF",  -- 175
        36745 => X"95",  -- 149
        36746 => X"A5",  -- 165
        36747 => X"9F",  -- 159
        36748 => X"99",  -- 153
        36749 => X"8F",  -- 143
        36750 => X"83",  -- 131
        36751 => X"8F",  -- 143
        36752 => X"88",  -- 136
        36753 => X"8B",  -- 139
        36754 => X"91",  -- 145
        36755 => X"8F",  -- 143
        36756 => X"83",  -- 131
        36757 => X"9B",  -- 155
        36758 => X"95",  -- 149
        36759 => X"91",  -- 145
        36760 => X"9D",  -- 157
        36761 => X"9E",  -- 158
        36762 => X"9C",  -- 156
        36763 => X"9B",  -- 155
        36764 => X"9C",  -- 156
        36765 => X"9F",  -- 159
        36766 => X"9D",  -- 157
        36767 => X"99",  -- 153
        36768 => X"A5",  -- 165
        36769 => X"A5",  -- 165
        36770 => X"AA",  -- 170
        36771 => X"A7",  -- 167
        36772 => X"A0",  -- 160
        36773 => X"AB",  -- 171
        36774 => X"B5",  -- 181
        36775 => X"B3",  -- 179
        36776 => X"9D",  -- 157
        36777 => X"9E",  -- 158
        36778 => X"8A",  -- 138
        36779 => X"7B",  -- 123
        36780 => X"71",  -- 113
        36781 => X"83",  -- 131
        36782 => X"A6",  -- 166
        36783 => X"AE",  -- 174
        36784 => X"C1",  -- 193
        36785 => X"C0",  -- 192
        36786 => X"C3",  -- 195
        36787 => X"C5",  -- 197
        36788 => X"C4",  -- 196
        36789 => X"C1",  -- 193
        36790 => X"C4",  -- 196
        36791 => X"C9",  -- 201
        36792 => X"D2",  -- 210
        36793 => X"CC",  -- 204
        36794 => X"C3",  -- 195
        36795 => X"BD",  -- 189
        36796 => X"AA",  -- 170
        36797 => X"80",  -- 128
        36798 => X"5E",  -- 94
        36799 => X"59",  -- 89
        36800 => X"5B",  -- 91
        36801 => X"5A",  -- 90
        36802 => X"59",  -- 89
        36803 => X"5B",  -- 91
        36804 => X"5D",  -- 93
        36805 => X"5F",  -- 95
        36806 => X"5E",  -- 94
        36807 => X"5D",  -- 93
        36808 => X"5B",  -- 91
        36809 => X"59",  -- 89
        36810 => X"57",  -- 87
        36811 => X"57",  -- 87
        36812 => X"59",  -- 89
        36813 => X"5A",  -- 90
        36814 => X"58",  -- 88
        36815 => X"56",  -- 86
        36816 => X"58",  -- 88
        36817 => X"57",  -- 87
        36818 => X"55",  -- 85
        36819 => X"57",  -- 87
        36820 => X"59",  -- 89
        36821 => X"57",  -- 87
        36822 => X"54",  -- 84
        36823 => X"50",  -- 80
        36824 => X"4E",  -- 78
        36825 => X"51",  -- 81
        36826 => X"62",  -- 98
        36827 => X"71",  -- 113
        36828 => X"7C",  -- 124
        36829 => X"87",  -- 135
        36830 => X"85",  -- 133
        36831 => X"75",  -- 117
        36832 => X"7F",  -- 127
        36833 => X"63",  -- 99
        36834 => X"41",  -- 65
        36835 => X"21",  -- 33
        36836 => X"18",  -- 24
        36837 => X"18",  -- 24
        36838 => X"2F",  -- 47
        36839 => X"69",  -- 105
        36840 => X"8D",  -- 141
        36841 => X"81",  -- 129
        36842 => X"5C",  -- 92
        36843 => X"23",  -- 35
        36844 => X"0E",  -- 14
        36845 => X"1B",  -- 27
        36846 => X"5F",  -- 95
        36847 => X"7E",  -- 126
        36848 => X"75",  -- 117
        36849 => X"6F",  -- 111
        36850 => X"47",  -- 71
        36851 => X"13",  -- 19
        36852 => X"03",  -- 3
        36853 => X"03",  -- 3
        36854 => X"0A",  -- 10
        36855 => X"20",  -- 32
        36856 => X"6F",  -- 111
        36857 => X"A2",  -- 162
        36858 => X"B1",  -- 177
        36859 => X"79",  -- 121
        36860 => X"33",  -- 51
        36861 => X"12",  -- 18
        36862 => X"11",  -- 17
        36863 => X"16",  -- 22
        36864 => X"31",  -- 49
        36865 => X"5C",  -- 92
        36866 => X"7B",  -- 123
        36867 => X"7D",  -- 125
        36868 => X"7F",  -- 127
        36869 => X"7C",  -- 124
        36870 => X"5A",  -- 90
        36871 => X"29",  -- 41
        36872 => X"13",  -- 19
        36873 => X"03",  -- 3
        36874 => X"24",  -- 36
        36875 => X"6C",  -- 108
        36876 => X"A3",  -- 163
        36877 => X"72",  -- 114
        36878 => X"41",  -- 65
        36879 => X"2D",  -- 45
        36880 => X"25",  -- 37
        36881 => X"2A",  -- 42
        36882 => X"26",  -- 38
        36883 => X"27",  -- 39
        36884 => X"35",  -- 53
        36885 => X"3F",  -- 63
        36886 => X"3F",  -- 63
        36887 => X"43",  -- 67
        36888 => X"59",  -- 89
        36889 => X"53",  -- 83
        36890 => X"4A",  -- 74
        36891 => X"5C",  -- 92
        36892 => X"58",  -- 88
        36893 => X"4B",  -- 75
        36894 => X"4E",  -- 78
        36895 => X"45",  -- 69
        36896 => X"41",  -- 65
        36897 => X"40",  -- 64
        36898 => X"46",  -- 70
        36899 => X"56",  -- 86
        36900 => X"46",  -- 70
        36901 => X"5D",  -- 93
        36902 => X"5E",  -- 94
        36903 => X"4F",  -- 79
        36904 => X"44",  -- 68
        36905 => X"4B",  -- 75
        36906 => X"4E",  -- 78
        36907 => X"42",  -- 66
        36908 => X"44",  -- 68
        36909 => X"46",  -- 70
        36910 => X"5E",  -- 94
        36911 => X"9F",  -- 159
        36912 => X"BC",  -- 188
        36913 => X"AF",  -- 175
        36914 => X"65",  -- 101
        36915 => X"08",  -- 8
        36916 => X"02",  -- 2
        36917 => X"0A",  -- 10
        36918 => X"28",  -- 40
        36919 => X"71",  -- 113
        36920 => X"AE",  -- 174
        36921 => X"B3",  -- 179
        36922 => X"A9",  -- 169
        36923 => X"A7",  -- 167
        36924 => X"9E",  -- 158
        36925 => X"6B",  -- 107
        36926 => X"2D",  -- 45
        36927 => X"0C",  -- 12
        36928 => X"16",  -- 22
        36929 => X"3C",  -- 60
        36930 => X"92",  -- 146
        36931 => X"CD",  -- 205
        36932 => X"DD",  -- 221
        36933 => X"A9",  -- 169
        36934 => X"3A",  -- 58
        36935 => X"00",  -- 0
        36936 => X"04",  -- 4
        36937 => X"06",  -- 6
        36938 => X"24",  -- 36
        36939 => X"8A",  -- 138
        36940 => X"C1",  -- 193
        36941 => X"BF",  -- 191
        36942 => X"CC",  -- 204
        36943 => X"C8",  -- 200
        36944 => X"C7",  -- 199
        36945 => X"9D",  -- 157
        36946 => X"3A",  -- 58
        36947 => X"1A",  -- 26
        36948 => X"2E",  -- 46
        36949 => X"93",  -- 147
        36950 => X"D1",  -- 209
        36951 => X"DE",  -- 222
        36952 => X"D4",  -- 212
        36953 => X"A5",  -- 165
        36954 => X"3A",  -- 58
        36955 => X"0B",  -- 11
        36956 => X"13",  -- 19
        36957 => X"16",  -- 22
        36958 => X"37",  -- 55
        36959 => X"6E",  -- 110
        36960 => X"96",  -- 150
        36961 => X"9F",  -- 159
        36962 => X"AE",  -- 174
        36963 => X"B9",  -- 185
        36964 => X"BD",  -- 189
        36965 => X"B8",  -- 184
        36966 => X"AF",  -- 175
        36967 => X"A9",  -- 169
        36968 => X"B3",  -- 179
        36969 => X"C4",  -- 196
        36970 => X"D2",  -- 210
        36971 => X"D0",  -- 208
        36972 => X"BC",  -- 188
        36973 => X"A5",  -- 165
        36974 => X"96",  -- 150
        36975 => X"90",  -- 144
        36976 => X"7B",  -- 123
        36977 => X"78",  -- 120
        36978 => X"6E",  -- 110
        36979 => X"5A",  -- 90
        36980 => X"41",  -- 65
        36981 => X"31",  -- 49
        36982 => X"34",  -- 52
        36983 => X"3E",  -- 62
        36984 => X"48",  -- 72
        36985 => X"52",  -- 82
        36986 => X"47",  -- 71
        36987 => X"43",  -- 67
        36988 => X"52",  -- 82
        36989 => X"3F",  -- 63
        36990 => X"29",  -- 41
        36991 => X"37",  -- 55
        36992 => X"25",  -- 37
        36993 => X"22",  -- 34
        36994 => X"26",  -- 38
        36995 => X"30",  -- 48
        36996 => X"35",  -- 53
        36997 => X"3D",  -- 61
        36998 => X"56",  -- 86
        36999 => X"72",  -- 114
        37000 => X"79",  -- 121
        37001 => X"8C",  -- 140
        37002 => X"92",  -- 146
        37003 => X"8C",  -- 140
        37004 => X"88",  -- 136
        37005 => X"87",  -- 135
        37006 => X"8D",  -- 141
        37007 => X"9A",  -- 154
        37008 => X"A4",  -- 164
        37009 => X"A1",  -- 161
        37010 => X"99",  -- 153
        37011 => X"93",  -- 147
        37012 => X"90",  -- 144
        37013 => X"90",  -- 144
        37014 => X"90",  -- 144
        37015 => X"8E",  -- 142
        37016 => X"A0",  -- 160
        37017 => X"99",  -- 153
        37018 => X"97",  -- 151
        37019 => X"9C",  -- 156
        37020 => X"9B",  -- 155
        37021 => X"8F",  -- 143
        37022 => X"81",  -- 129
        37023 => X"79",  -- 121
        37024 => X"70",  -- 112
        37025 => X"74",  -- 116
        37026 => X"76",  -- 118
        37027 => X"72",  -- 114
        37028 => X"69",  -- 105
        37029 => X"60",  -- 96
        37030 => X"5A",  -- 90
        37031 => X"58",  -- 88
        37032 => X"53",  -- 83
        37033 => X"54",  -- 84
        37034 => X"4E",  -- 78
        37035 => X"3F",  -- 63
        37036 => X"32",  -- 50
        37037 => X"34",  -- 52
        37038 => X"45",  -- 69
        37039 => X"54",  -- 84
        37040 => X"67",  -- 103
        37041 => X"7E",  -- 126
        37042 => X"8C",  -- 140
        37043 => X"9A",  -- 154
        37044 => X"9C",  -- 156
        37045 => X"9E",  -- 158
        37046 => X"AE",  -- 174
        37047 => X"B2",  -- 178
        37048 => X"B4",  -- 180
        37049 => X"BC",  -- 188
        37050 => X"B9",  -- 185
        37051 => X"BD",  -- 189
        37052 => X"B7",  -- 183
        37053 => X"C2",  -- 194
        37054 => X"BA",  -- 186
        37055 => X"B5",  -- 181
        37056 => X"B1",  -- 177
        37057 => X"B0",  -- 176
        37058 => X"BC",  -- 188
        37059 => X"B5",  -- 181
        37060 => X"B5",  -- 181
        37061 => X"A1",  -- 161
        37062 => X"A9",  -- 169
        37063 => X"AF",  -- 175
        37064 => X"A7",  -- 167
        37065 => X"93",  -- 147
        37066 => X"A7",  -- 167
        37067 => X"9E",  -- 158
        37068 => X"9B",  -- 155
        37069 => X"8D",  -- 141
        37070 => X"8E",  -- 142
        37071 => X"93",  -- 147
        37072 => X"8A",  -- 138
        37073 => X"8E",  -- 142
        37074 => X"96",  -- 150
        37075 => X"95",  -- 149
        37076 => X"88",  -- 136
        37077 => X"9F",  -- 159
        37078 => X"9B",  -- 155
        37079 => X"9D",  -- 157
        37080 => X"9E",  -- 158
        37081 => X"A2",  -- 162
        37082 => X"A1",  -- 161
        37083 => X"98",  -- 152
        37084 => X"9D",  -- 157
        37085 => X"A8",  -- 168
        37086 => X"A6",  -- 166
        37087 => X"99",  -- 153
        37088 => X"A7",  -- 167
        37089 => X"AC",  -- 172
        37090 => X"B0",  -- 176
        37091 => X"AD",  -- 173
        37092 => X"A8",  -- 168
        37093 => X"B0",  -- 176
        37094 => X"BC",  -- 188
        37095 => X"BE",  -- 190
        37096 => X"A3",  -- 163
        37097 => X"99",  -- 153
        37098 => X"8E",  -- 142
        37099 => X"7D",  -- 125
        37100 => X"67",  -- 103
        37101 => X"75",  -- 117
        37102 => X"9A",  -- 154
        37103 => X"A8",  -- 168
        37104 => X"BD",  -- 189
        37105 => X"C3",  -- 195
        37106 => X"CC",  -- 204
        37107 => X"CD",  -- 205
        37108 => X"C3",  -- 195
        37109 => X"B8",  -- 184
        37110 => X"BF",  -- 191
        37111 => X"CE",  -- 206
        37112 => X"CC",  -- 204
        37113 => X"C8",  -- 200
        37114 => X"BF",  -- 191
        37115 => X"B4",  -- 180
        37116 => X"A1",  -- 161
        37117 => X"84",  -- 132
        37118 => X"67",  -- 103
        37119 => X"59",  -- 89
        37120 => X"5F",  -- 95
        37121 => X"5E",  -- 94
        37122 => X"5E",  -- 94
        37123 => X"5E",  -- 94
        37124 => X"5E",  -- 94
        37125 => X"5C",  -- 92
        37126 => X"5A",  -- 90
        37127 => X"58",  -- 88
        37128 => X"5B",  -- 91
        37129 => X"59",  -- 89
        37130 => X"57",  -- 87
        37131 => X"57",  -- 87
        37132 => X"59",  -- 89
        37133 => X"59",  -- 89
        37134 => X"57",  -- 87
        37135 => X"54",  -- 84
        37136 => X"54",  -- 84
        37137 => X"53",  -- 83
        37138 => X"52",  -- 82
        37139 => X"54",  -- 84
        37140 => X"58",  -- 88
        37141 => X"57",  -- 87
        37142 => X"55",  -- 85
        37143 => X"51",  -- 81
        37144 => X"53",  -- 83
        37145 => X"4F",  -- 79
        37146 => X"5B",  -- 91
        37147 => X"6F",  -- 111
        37148 => X"79",  -- 121
        37149 => X"81",  -- 129
        37150 => X"87",  -- 135
        37151 => X"85",  -- 133
        37152 => X"7D",  -- 125
        37153 => X"65",  -- 101
        37154 => X"46",  -- 70
        37155 => X"25",  -- 37
        37156 => X"16",  -- 22
        37157 => X"14",  -- 20
        37158 => X"2E",  -- 46
        37159 => X"6E",  -- 110
        37160 => X"95",  -- 149
        37161 => X"8B",  -- 139
        37162 => X"69",  -- 105
        37163 => X"2A",  -- 42
        37164 => X"0D",  -- 13
        37165 => X"1E",  -- 30
        37166 => X"60",  -- 96
        37167 => X"72",  -- 114
        37168 => X"7C",  -- 124
        37169 => X"7A",  -- 122
        37170 => X"4C",  -- 76
        37171 => X"1C",  -- 28
        37172 => X"0F",  -- 15
        37173 => X"0E",  -- 14
        37174 => X"13",  -- 19
        37175 => X"1B",  -- 27
        37176 => X"3C",  -- 60
        37177 => X"94",  -- 148
        37178 => X"B7",  -- 183
        37179 => X"9D",  -- 157
        37180 => X"75",  -- 117
        37181 => X"2C",  -- 44
        37182 => X"01",  -- 1
        37183 => X"16",  -- 22
        37184 => X"0F",  -- 15
        37185 => X"1C",  -- 28
        37186 => X"37",  -- 55
        37187 => X"53",  -- 83
        37188 => X"54",  -- 84
        37189 => X"38",  -- 56
        37190 => X"1C",  -- 28
        37191 => X"0C",  -- 12
        37192 => X"0D",  -- 13
        37193 => X"01",  -- 1
        37194 => X"10",  -- 16
        37195 => X"54",  -- 84
        37196 => X"A4",  -- 164
        37197 => X"86",  -- 134
        37198 => X"4B",  -- 75
        37199 => X"2E",  -- 46
        37200 => X"27",  -- 39
        37201 => X"27",  -- 39
        37202 => X"2B",  -- 43
        37203 => X"35",  -- 53
        37204 => X"3F",  -- 63
        37205 => X"3A",  -- 58
        37206 => X"37",  -- 55
        37207 => X"44",  -- 68
        37208 => X"5A",  -- 90
        37209 => X"44",  -- 68
        37210 => X"52",  -- 82
        37211 => X"57",  -- 87
        37212 => X"56",  -- 86
        37213 => X"51",  -- 81
        37214 => X"46",  -- 70
        37215 => X"48",  -- 72
        37216 => X"45",  -- 69
        37217 => X"40",  -- 64
        37218 => X"42",  -- 66
        37219 => X"53",  -- 83
        37220 => X"48",  -- 72
        37221 => X"62",  -- 98
        37222 => X"63",  -- 99
        37223 => X"52",  -- 82
        37224 => X"5A",  -- 90
        37225 => X"59",  -- 89
        37226 => X"4E",  -- 78
        37227 => X"3E",  -- 62
        37228 => X"42",  -- 66
        37229 => X"55",  -- 85
        37230 => X"79",  -- 121
        37231 => X"C1",  -- 193
        37232 => X"CD",  -- 205
        37233 => X"C2",  -- 194
        37234 => X"52",  -- 82
        37235 => X"0C",  -- 12
        37236 => X"14",  -- 20
        37237 => X"08",  -- 8
        37238 => X"04",  -- 4
        37239 => X"1D",  -- 29
        37240 => X"42",  -- 66
        37241 => X"74",  -- 116
        37242 => X"8B",  -- 139
        37243 => X"6B",  -- 107
        37244 => X"40",  -- 64
        37245 => X"1C",  -- 28
        37246 => X"10",  -- 16
        37247 => X"21",  -- 33
        37248 => X"2C",  -- 44
        37249 => X"6F",  -- 111
        37250 => X"C5",  -- 197
        37251 => X"D3",  -- 211
        37252 => X"B5",  -- 181
        37253 => X"77",  -- 119
        37254 => X"26",  -- 38
        37255 => X"0E",  -- 14
        37256 => X"0F",  -- 15
        37257 => X"05",  -- 5
        37258 => X"29",  -- 41
        37259 => X"8D",  -- 141
        37260 => X"C0",  -- 192
        37261 => X"BF",  -- 191
        37262 => X"C1",  -- 193
        37263 => X"AD",  -- 173
        37264 => X"C7",  -- 199
        37265 => X"9F",  -- 159
        37266 => X"3B",  -- 59
        37267 => X"29",  -- 41
        37268 => X"41",  -- 65
        37269 => X"A3",  -- 163
        37270 => X"D1",  -- 209
        37271 => X"E0",  -- 224
        37272 => X"DA",  -- 218
        37273 => X"B8",  -- 184
        37274 => X"53",  -- 83
        37275 => X"0D",  -- 13
        37276 => X"16",  -- 22
        37277 => X"1B",  -- 27
        37278 => X"37",  -- 55
        37279 => X"6A",  -- 106
        37280 => X"96",  -- 150
        37281 => X"A5",  -- 165
        37282 => X"B6",  -- 182
        37283 => X"BD",  -- 189
        37284 => X"C0",  -- 192
        37285 => X"C0",  -- 192
        37286 => X"B3",  -- 179
        37287 => X"A6",  -- 166
        37288 => X"AC",  -- 172
        37289 => X"BD",  -- 189
        37290 => X"CF",  -- 207
        37291 => X"CF",  -- 207
        37292 => X"BF",  -- 191
        37293 => X"A7",  -- 167
        37294 => X"94",  -- 148
        37295 => X"89",  -- 137
        37296 => X"8E",  -- 142
        37297 => X"7C",  -- 124
        37298 => X"64",  -- 100
        37299 => X"4E",  -- 78
        37300 => X"3C",  -- 60
        37301 => X"32",  -- 50
        37302 => X"33",  -- 51
        37303 => X"38",  -- 56
        37304 => X"4A",  -- 74
        37305 => X"5A",  -- 90
        37306 => X"49",  -- 73
        37307 => X"3C",  -- 60
        37308 => X"53",  -- 83
        37309 => X"50",  -- 80
        37310 => X"2F",  -- 47
        37311 => X"23",  -- 35
        37312 => X"29",  -- 41
        37313 => X"24",  -- 36
        37314 => X"28",  -- 40
        37315 => X"36",  -- 54
        37316 => X"41",  -- 65
        37317 => X"4C",  -- 76
        37318 => X"60",  -- 96
        37319 => X"75",  -- 117
        37320 => X"7D",  -- 125
        37321 => X"8E",  -- 142
        37322 => X"93",  -- 147
        37323 => X"8D",  -- 141
        37324 => X"88",  -- 136
        37325 => X"83",  -- 131
        37326 => X"86",  -- 134
        37327 => X"91",  -- 145
        37328 => X"9C",  -- 156
        37329 => X"A0",  -- 160
        37330 => X"9B",  -- 155
        37331 => X"8F",  -- 143
        37332 => X"8F",  -- 143
        37333 => X"95",  -- 149
        37334 => X"91",  -- 145
        37335 => X"84",  -- 132
        37336 => X"92",  -- 146
        37337 => X"95",  -- 149
        37338 => X"93",  -- 147
        37339 => X"8D",  -- 141
        37340 => X"89",  -- 137
        37341 => X"85",  -- 133
        37342 => X"7A",  -- 122
        37343 => X"6E",  -- 110
        37344 => X"65",  -- 101
        37345 => X"67",  -- 103
        37346 => X"69",  -- 105
        37347 => X"6A",  -- 106
        37348 => X"67",  -- 103
        37349 => X"5F",  -- 95
        37350 => X"57",  -- 87
        37351 => X"52",  -- 82
        37352 => X"4C",  -- 76
        37353 => X"4A",  -- 74
        37354 => X"42",  -- 66
        37355 => X"36",  -- 54
        37356 => X"2A",  -- 42
        37357 => X"30",  -- 48
        37358 => X"45",  -- 69
        37359 => X"59",  -- 89
        37360 => X"70",  -- 112
        37361 => X"88",  -- 136
        37362 => X"93",  -- 147
        37363 => X"9F",  -- 159
        37364 => X"A3",  -- 163
        37365 => X"A6",  -- 166
        37366 => X"B3",  -- 179
        37367 => X"B3",  -- 179
        37368 => X"B5",  -- 181
        37369 => X"C2",  -- 194
        37370 => X"BB",  -- 187
        37371 => X"C2",  -- 194
        37372 => X"B2",  -- 178
        37373 => X"BF",  -- 191
        37374 => X"B4",  -- 180
        37375 => X"B3",  -- 179
        37376 => X"B1",  -- 177
        37377 => X"A9",  -- 169
        37378 => X"B4",  -- 180
        37379 => X"B0",  -- 176
        37380 => X"B7",  -- 183
        37381 => X"A3",  -- 163
        37382 => X"A4",  -- 164
        37383 => X"A4",  -- 164
        37384 => X"9F",  -- 159
        37385 => X"96",  -- 150
        37386 => X"A8",  -- 168
        37387 => X"9E",  -- 158
        37388 => X"9C",  -- 156
        37389 => X"90",  -- 144
        37390 => X"96",  -- 150
        37391 => X"96",  -- 150
        37392 => X"8D",  -- 141
        37393 => X"8F",  -- 143
        37394 => X"96",  -- 150
        37395 => X"98",  -- 152
        37396 => X"8A",  -- 138
        37397 => X"9F",  -- 159
        37398 => X"9D",  -- 157
        37399 => X"A3",  -- 163
        37400 => X"AB",  -- 171
        37401 => X"9C",  -- 156
        37402 => X"98",  -- 152
        37403 => X"A4",  -- 164
        37404 => X"A9",  -- 169
        37405 => X"A4",  -- 164
        37406 => X"9F",  -- 159
        37407 => X"A5",  -- 165
        37408 => X"A3",  -- 163
        37409 => X"AC",  -- 172
        37410 => X"B2",  -- 178
        37411 => X"B0",  -- 176
        37412 => X"B2",  -- 178
        37413 => X"B7",  -- 183
        37414 => X"BD",  -- 189
        37415 => X"C3",  -- 195
        37416 => X"B7",  -- 183
        37417 => X"9D",  -- 157
        37418 => X"93",  -- 147
        37419 => X"81",  -- 129
        37420 => X"69",  -- 105
        37421 => X"6F",  -- 111
        37422 => X"8F",  -- 143
        37423 => X"A9",  -- 169
        37424 => X"B8",  -- 184
        37425 => X"C0",  -- 192
        37426 => X"CB",  -- 203
        37427 => X"CE",  -- 206
        37428 => X"C1",  -- 193
        37429 => X"B5",  -- 181
        37430 => X"B9",  -- 185
        37431 => X"C6",  -- 198
        37432 => X"C4",  -- 196
        37433 => X"C7",  -- 199
        37434 => X"C0",  -- 192
        37435 => X"AA",  -- 170
        37436 => X"92",  -- 146
        37437 => X"84",  -- 132
        37438 => X"72",  -- 114
        37439 => X"5F",  -- 95
        37440 => X"5B",  -- 91
        37441 => X"5B",  -- 91
        37442 => X"5B",  -- 91
        37443 => X"5B",  -- 91
        37444 => X"59",  -- 89
        37445 => X"57",  -- 87
        37446 => X"55",  -- 85
        37447 => X"54",  -- 84
        37448 => X"57",  -- 87
        37449 => X"57",  -- 87
        37450 => X"58",  -- 88
        37451 => X"59",  -- 89
        37452 => X"5A",  -- 90
        37453 => X"5A",  -- 90
        37454 => X"57",  -- 87
        37455 => X"56",  -- 86
        37456 => X"51",  -- 81
        37457 => X"50",  -- 80
        37458 => X"4F",  -- 79
        37459 => X"51",  -- 81
        37460 => X"54",  -- 84
        37461 => X"54",  -- 84
        37462 => X"51",  -- 81
        37463 => X"4E",  -- 78
        37464 => X"50",  -- 80
        37465 => X"47",  -- 71
        37466 => X"55",  -- 85
        37467 => X"70",  -- 112
        37468 => X"7B",  -- 123
        37469 => X"7E",  -- 126
        37470 => X"86",  -- 134
        37471 => X"8C",  -- 140
        37472 => X"76",  -- 118
        37473 => X"6D",  -- 109
        37474 => X"50",  -- 80
        37475 => X"21",  -- 33
        37476 => X"0F",  -- 15
        37477 => X"18",  -- 24
        37478 => X"33",  -- 51
        37479 => X"67",  -- 103
        37480 => X"94",  -- 148
        37481 => X"8F",  -- 143
        37482 => X"67",  -- 103
        37483 => X"21",  -- 33
        37484 => X"08",  -- 8
        37485 => X"20",  -- 32
        37486 => X"64",  -- 100
        37487 => X"75",  -- 117
        37488 => X"75",  -- 117
        37489 => X"6E",  -- 110
        37490 => X"35",  -- 53
        37491 => X"09",  -- 9
        37492 => X"05",  -- 5
        37493 => X"0B",  -- 11
        37494 => X"10",  -- 16
        37495 => X"0E",  -- 14
        37496 => X"0B",  -- 11
        37497 => X"4B",  -- 75
        37498 => X"96",  -- 150
        37499 => X"BE",  -- 190
        37500 => X"A4",  -- 164
        37501 => X"58",  -- 88
        37502 => X"1B",  -- 27
        37503 => X"10",  -- 16
        37504 => X"0E",  -- 14
        37505 => X"07",  -- 7
        37506 => X"04",  -- 4
        37507 => X"09",  -- 9
        37508 => X"0A",  -- 10
        37509 => X"05",  -- 5
        37510 => X"04",  -- 4
        37511 => X"09",  -- 9
        37512 => X"06",  -- 6
        37513 => X"02",  -- 2
        37514 => X"0C",  -- 12
        37515 => X"45",  -- 69
        37516 => X"A4",  -- 164
        37517 => X"95",  -- 149
        37518 => X"54",  -- 84
        37519 => X"31",  -- 49
        37520 => X"29",  -- 41
        37521 => X"28",  -- 40
        37522 => X"29",  -- 41
        37523 => X"35",  -- 53
        37524 => X"3A",  -- 58
        37525 => X"30",  -- 48
        37526 => X"32",  -- 50
        37527 => X"47",  -- 71
        37528 => X"54",  -- 84
        37529 => X"3D",  -- 61
        37530 => X"55",  -- 85
        37531 => X"50",  -- 80
        37532 => X"53",  -- 83
        37533 => X"4F",  -- 79
        37534 => X"44",  -- 68
        37535 => X"4B",  -- 75
        37536 => X"59",  -- 89
        37537 => X"50",  -- 80
        37538 => X"51",  -- 81
        37539 => X"58",  -- 88
        37540 => X"50",  -- 80
        37541 => X"5D",  -- 93
        37542 => X"5C",  -- 92
        37543 => X"4E",  -- 78
        37544 => X"5F",  -- 95
        37545 => X"57",  -- 87
        37546 => X"46",  -- 70
        37547 => X"3B",  -- 59
        37548 => X"3F",  -- 63
        37549 => X"61",  -- 97
        37550 => X"8A",  -- 138
        37551 => X"D0",  -- 208
        37552 => X"DA",  -- 218
        37553 => X"C1",  -- 193
        37554 => X"3B",  -- 59
        37555 => X"13",  -- 19
        37556 => X"15",  -- 21
        37557 => X"08",  -- 8
        37558 => X"05",  -- 5
        37559 => X"0B",  -- 11
        37560 => X"0D",  -- 13
        37561 => X"0C",  -- 12
        37562 => X"0D",  -- 13
        37563 => X"0C",  -- 12
        37564 => X"18",  -- 24
        37565 => X"1C",  -- 28
        37566 => X"1E",  -- 30
        37567 => X"3B",  -- 59
        37568 => X"84",  -- 132
        37569 => X"B4",  -- 180
        37570 => X"E8",  -- 232
        37571 => X"B9",  -- 185
        37572 => X"53",  -- 83
        37573 => X"1A",  -- 26
        37574 => X"0B",  -- 11
        37575 => X"0A",  -- 10
        37576 => X"02",  -- 2
        37577 => X"15",  -- 21
        37578 => X"4A",  -- 74
        37579 => X"8F",  -- 143
        37580 => X"B3",  -- 179
        37581 => X"C1",  -- 193
        37582 => X"C8",  -- 200
        37583 => X"B4",  -- 180
        37584 => X"B9",  -- 185
        37585 => X"94",  -- 148
        37586 => X"2B",  -- 43
        37587 => X"1F",  -- 31
        37588 => X"40",  -- 64
        37589 => X"A7",  -- 167
        37590 => X"CC",  -- 204
        37591 => X"D9",  -- 217
        37592 => X"DE",  -- 222
        37593 => X"CD",  -- 205
        37594 => X"76",  -- 118
        37595 => X"19",  -- 25
        37596 => X"1A",  -- 26
        37597 => X"26",  -- 38
        37598 => X"46",  -- 70
        37599 => X"6F",  -- 111
        37600 => X"93",  -- 147
        37601 => X"A6",  -- 166
        37602 => X"B9",  -- 185
        37603 => X"C0",  -- 192
        37604 => X"C3",  -- 195
        37605 => X"C6",  -- 198
        37606 => X"BA",  -- 186
        37607 => X"AA",  -- 170
        37608 => X"AB",  -- 171
        37609 => X"B9",  -- 185
        37610 => X"C9",  -- 201
        37611 => X"CF",  -- 207
        37612 => X"C6",  -- 198
        37613 => X"AF",  -- 175
        37614 => X"97",  -- 151
        37615 => X"87",  -- 135
        37616 => X"84",  -- 132
        37617 => X"77",  -- 119
        37618 => X"63",  -- 99
        37619 => X"4F",  -- 79
        37620 => X"3F",  -- 63
        37621 => X"38",  -- 56
        37622 => X"3F",  -- 63
        37623 => X"48",  -- 72
        37624 => X"49",  -- 73
        37625 => X"4C",  -- 76
        37626 => X"58",  -- 88
        37627 => X"4B",  -- 75
        37628 => X"38",  -- 56
        37629 => X"44",  -- 68
        37630 => X"48",  -- 72
        37631 => X"2A",  -- 42
        37632 => X"26",  -- 38
        37633 => X"25",  -- 37
        37634 => X"2A",  -- 42
        37635 => X"38",  -- 56
        37636 => X"4C",  -- 76
        37637 => X"5D",  -- 93
        37638 => X"6A",  -- 106
        37639 => X"75",  -- 117
        37640 => X"80",  -- 128
        37641 => X"8E",  -- 142
        37642 => X"91",  -- 145
        37643 => X"8E",  -- 142
        37644 => X"8A",  -- 138
        37645 => X"82",  -- 130
        37646 => X"81",  -- 129
        37647 => X"8A",  -- 138
        37648 => X"88",  -- 136
        37649 => X"98",  -- 152
        37650 => X"9E",  -- 158
        37651 => X"94",  -- 148
        37652 => X"8C",  -- 140
        37653 => X"8F",  -- 143
        37654 => X"8F",  -- 143
        37655 => X"88",  -- 136
        37656 => X"87",  -- 135
        37657 => X"8A",  -- 138
        37658 => X"84",  -- 132
        37659 => X"76",  -- 118
        37660 => X"72",  -- 114
        37661 => X"76",  -- 118
        37662 => X"75",  -- 117
        37663 => X"6D",  -- 109
        37664 => X"69",  -- 105
        37665 => X"64",  -- 100
        37666 => X"5F",  -- 95
        37667 => X"60",  -- 96
        37668 => X"5F",  -- 95
        37669 => X"5A",  -- 90
        37670 => X"54",  -- 84
        37671 => X"51",  -- 81
        37672 => X"44",  -- 68
        37673 => X"41",  -- 65
        37674 => X"3A",  -- 58
        37675 => X"33",  -- 51
        37676 => X"2F",  -- 47
        37677 => X"34",  -- 52
        37678 => X"45",  -- 69
        37679 => X"54",  -- 84
        37680 => X"6D",  -- 109
        37681 => X"87",  -- 135
        37682 => X"98",  -- 152
        37683 => X"A9",  -- 169
        37684 => X"AF",  -- 175
        37685 => X"B0",  -- 176
        37686 => X"B9",  -- 185
        37687 => X"B3",  -- 179
        37688 => X"BE",  -- 190
        37689 => X"C4",  -- 196
        37690 => X"BC",  -- 188
        37691 => X"C0",  -- 192
        37692 => X"B1",  -- 177
        37693 => X"BB",  -- 187
        37694 => X"B5",  -- 181
        37695 => X"B9",  -- 185
        37696 => X"AF",  -- 175
        37697 => X"A5",  -- 165
        37698 => X"A5",  -- 165
        37699 => X"AB",  -- 171
        37700 => X"B1",  -- 177
        37701 => X"A4",  -- 164
        37702 => X"9E",  -- 158
        37703 => X"9D",  -- 157
        37704 => X"9A",  -- 154
        37705 => X"9A",  -- 154
        37706 => X"A4",  -- 164
        37707 => X"A1",  -- 161
        37708 => X"9A",  -- 154
        37709 => X"96",  -- 150
        37710 => X"9B",  -- 155
        37711 => X"95",  -- 149
        37712 => X"95",  -- 149
        37713 => X"91",  -- 145
        37714 => X"96",  -- 150
        37715 => X"99",  -- 153
        37716 => X"8B",  -- 139
        37717 => X"9D",  -- 157
        37718 => X"9B",  -- 155
        37719 => X"A3",  -- 163
        37720 => X"A9",  -- 169
        37721 => X"A1",  -- 161
        37722 => X"9D",  -- 157
        37723 => X"A0",  -- 160
        37724 => X"A6",  -- 166
        37725 => X"A7",  -- 167
        37726 => X"A5",  -- 165
        37727 => X"A4",  -- 164
        37728 => X"A2",  -- 162
        37729 => X"AB",  -- 171
        37730 => X"AD",  -- 173
        37731 => X"B0",  -- 176
        37732 => X"B9",  -- 185
        37733 => X"BC",  -- 188
        37734 => X"BB",  -- 187
        37735 => X"C0",  -- 192
        37736 => X"B7",  -- 183
        37737 => X"9B",  -- 155
        37738 => X"95",  -- 149
        37739 => X"8D",  -- 141
        37740 => X"7E",  -- 126
        37741 => X"7B",  -- 123
        37742 => X"84",  -- 132
        37743 => X"9C",  -- 156
        37744 => X"BB",  -- 187
        37745 => X"BE",  -- 190
        37746 => X"C3",  -- 195
        37747 => X"C7",  -- 199
        37748 => X"C3",  -- 195
        37749 => X"BB",  -- 187
        37750 => X"B8",  -- 184
        37751 => X"B9",  -- 185
        37752 => X"BF",  -- 191
        37753 => X"C4",  -- 196
        37754 => X"C2",  -- 194
        37755 => X"A6",  -- 166
        37756 => X"85",  -- 133
        37757 => X"79",  -- 121
        37758 => X"73",  -- 115
        37759 => X"66",  -- 102
        37760 => X"50",  -- 80
        37761 => X"51",  -- 81
        37762 => X"53",  -- 83
        37763 => X"53",  -- 83
        37764 => X"53",  -- 83
        37765 => X"52",  -- 82
        37766 => X"51",  -- 81
        37767 => X"52",  -- 82
        37768 => X"52",  -- 82
        37769 => X"55",  -- 85
        37770 => X"58",  -- 88
        37771 => X"59",  -- 89
        37772 => X"58",  -- 88
        37773 => X"56",  -- 86
        37774 => X"55",  -- 85
        37775 => X"53",  -- 83
        37776 => X"4B",  -- 75
        37777 => X"4B",  -- 75
        37778 => X"4C",  -- 76
        37779 => X"4E",  -- 78
        37780 => X"53",  -- 83
        37781 => X"53",  -- 83
        37782 => X"51",  -- 81
        37783 => X"4E",  -- 78
        37784 => X"4C",  -- 76
        37785 => X"45",  -- 69
        37786 => X"54",  -- 84
        37787 => X"6D",  -- 109
        37788 => X"77",  -- 119
        37789 => X"7B",  -- 123
        37790 => X"83",  -- 131
        37791 => X"8A",  -- 138
        37792 => X"76",  -- 118
        37793 => X"6D",  -- 109
        37794 => X"4F",  -- 79
        37795 => X"21",  -- 33
        37796 => X"0F",  -- 15
        37797 => X"17",  -- 23
        37798 => X"2F",  -- 47
        37799 => X"61",  -- 97
        37800 => X"8A",  -- 138
        37801 => X"8E",  -- 142
        37802 => X"64",  -- 100
        37803 => X"1B",  -- 27
        37804 => X"08",  -- 8
        37805 => X"26",  -- 38
        37806 => X"6A",  -- 106
        37807 => X"7C",  -- 124
        37808 => X"6F",  -- 111
        37809 => X"64",  -- 100
        37810 => X"26",  -- 38
        37811 => X"07",  -- 7
        37812 => X"17",  -- 23
        37813 => X"30",  -- 48
        37814 => X"42",  -- 66
        37815 => X"3D",  -- 61
        37816 => X"16",  -- 22
        37817 => X"11",  -- 17
        37818 => X"5C",  -- 92
        37819 => X"AE",  -- 174
        37820 => X"AE",  -- 174
        37821 => X"8F",  -- 143
        37822 => X"6A",  -- 106
        37823 => X"3A",  -- 58
        37824 => X"20",  -- 32
        37825 => X"20",  -- 32
        37826 => X"17",  -- 23
        37827 => X"0F",  -- 15
        37828 => X"11",  -- 17
        37829 => X"19",  -- 25
        37830 => X"12",  -- 18
        37831 => X"05",  -- 5
        37832 => X"0D",  -- 13
        37833 => X"0B",  -- 11
        37834 => X"0A",  -- 10
        37835 => X"37",  -- 55
        37836 => X"98",  -- 152
        37837 => X"8E",  -- 142
        37838 => X"52",  -- 82
        37839 => X"35",  -- 53
        37840 => X"2A",  -- 42
        37841 => X"29",  -- 41
        37842 => X"27",  -- 39
        37843 => X"2D",  -- 45
        37844 => X"32",  -- 50
        37845 => X"2E",  -- 46
        37846 => X"34",  -- 52
        37847 => X"45",  -- 69
        37848 => X"4D",  -- 77
        37849 => X"43",  -- 67
        37850 => X"52",  -- 82
        37851 => X"4C",  -- 76
        37852 => X"4D",  -- 77
        37853 => X"45",  -- 69
        37854 => X"4F",  -- 79
        37855 => X"4F",  -- 79
        37856 => X"5A",  -- 90
        37857 => X"56",  -- 86
        37858 => X"5C",  -- 92
        37859 => X"5B",  -- 91
        37860 => X"5B",  -- 91
        37861 => X"52",  -- 82
        37862 => X"51",  -- 81
        37863 => X"4B",  -- 75
        37864 => X"53",  -- 83
        37865 => X"49",  -- 73
        37866 => X"42",  -- 66
        37867 => X"43",  -- 67
        37868 => X"3F",  -- 63
        37869 => X"67",  -- 103
        37870 => X"90",  -- 144
        37871 => X"C9",  -- 201
        37872 => X"D7",  -- 215
        37873 => X"9D",  -- 157
        37874 => X"18",  -- 24
        37875 => X"19",  -- 25
        37876 => X"12",  -- 18
        37877 => X"16",  -- 22
        37878 => X"17",  -- 23
        37879 => X"1E",  -- 30
        37880 => X"12",  -- 18
        37881 => X"0D",  -- 13
        37882 => X"1D",  -- 29
        37883 => X"1F",  -- 31
        37884 => X"1D",  -- 29
        37885 => X"28",  -- 40
        37886 => X"4D",  -- 77
        37887 => X"90",  -- 144
        37888 => X"B5",  -- 181
        37889 => X"CE",  -- 206
        37890 => X"BA",  -- 186
        37891 => X"74",  -- 116
        37892 => X"2A",  -- 42
        37893 => X"09",  -- 9
        37894 => X"10",  -- 16
        37895 => X"10",  -- 16
        37896 => X"13",  -- 19
        37897 => X"3B",  -- 59
        37898 => X"85",  -- 133
        37899 => X"B1",  -- 177
        37900 => X"BD",  -- 189
        37901 => X"C5",  -- 197
        37902 => X"BE",  -- 190
        37903 => X"BA",  -- 186
        37904 => X"B4",  -- 180
        37905 => X"95",  -- 149
        37906 => X"22",  -- 34
        37907 => X"0F",  -- 15
        37908 => X"32",  -- 50
        37909 => X"A9",  -- 169
        37910 => X"CD",  -- 205
        37911 => X"D3",  -- 211
        37912 => X"D9",  -- 217
        37913 => X"D8",  -- 216
        37914 => X"93",  -- 147
        37915 => X"24",  -- 36
        37916 => X"17",  -- 23
        37917 => X"2C",  -- 44
        37918 => X"56",  -- 86
        37919 => X"7D",  -- 125
        37920 => X"9A",  -- 154
        37921 => X"A6",  -- 166
        37922 => X"B7",  -- 183
        37923 => X"C0",  -- 192
        37924 => X"C4",  -- 196
        37925 => X"BF",  -- 191
        37926 => X"B7",  -- 183
        37927 => X"B2",  -- 178
        37928 => X"B2",  -- 178
        37929 => X"BA",  -- 186
        37930 => X"C7",  -- 199
        37931 => X"D0",  -- 208
        37932 => X"CE",  -- 206
        37933 => X"B8",  -- 184
        37934 => X"9C",  -- 156
        37935 => X"86",  -- 134
        37936 => X"70",  -- 112
        37937 => X"6A",  -- 106
        37938 => X"62",  -- 98
        37939 => X"55",  -- 85
        37940 => X"48",  -- 72
        37941 => X"44",  -- 68
        37942 => X"4E",  -- 78
        37943 => X"5C",  -- 92
        37944 => X"50",  -- 80
        37945 => X"44",  -- 68
        37946 => X"58",  -- 88
        37947 => X"55",  -- 85
        37948 => X"33",  -- 51
        37949 => X"37",  -- 55
        37950 => X"49",  -- 73
        37951 => X"3B",  -- 59
        37952 => X"29",  -- 41
        37953 => X"2E",  -- 46
        37954 => X"34",  -- 52
        37955 => X"40",  -- 64
        37956 => X"52",  -- 82
        37957 => X"65",  -- 101
        37958 => X"6D",  -- 109
        37959 => X"70",  -- 112
        37960 => X"7D",  -- 125
        37961 => X"88",  -- 136
        37962 => X"8A",  -- 138
        37963 => X"89",  -- 137
        37964 => X"87",  -- 135
        37965 => X"7F",  -- 127
        37966 => X"7C",  -- 124
        37967 => X"83",  -- 131
        37968 => X"7E",  -- 126
        37969 => X"8A",  -- 138
        37970 => X"95",  -- 149
        37971 => X"94",  -- 148
        37972 => X"8B",  -- 139
        37973 => X"82",  -- 130
        37974 => X"84",  -- 132
        37975 => X"8A",  -- 138
        37976 => X"83",  -- 131
        37977 => X"7E",  -- 126
        37978 => X"74",  -- 116
        37979 => X"6B",  -- 107
        37980 => X"68",  -- 104
        37981 => X"69",  -- 105
        37982 => X"6A",  -- 106
        37983 => X"6A",  -- 106
        37984 => X"67",  -- 103
        37985 => X"60",  -- 96
        37986 => X"5D",  -- 93
        37987 => X"5E",  -- 94
        37988 => X"5B",  -- 91
        37989 => X"55",  -- 85
        37990 => X"51",  -- 81
        37991 => X"4E",  -- 78
        37992 => X"43",  -- 67
        37993 => X"3D",  -- 61
        37994 => X"38",  -- 56
        37995 => X"3B",  -- 59
        37996 => X"3E",  -- 62
        37997 => X"40",  -- 64
        37998 => X"45",  -- 69
        37999 => X"4B",  -- 75
        38000 => X"65",  -- 101
        38001 => X"87",  -- 135
        38002 => X"9D",  -- 157
        38003 => X"AD",  -- 173
        38004 => X"B1",  -- 177
        38005 => X"B2",  -- 178
        38006 => X"BD",  -- 189
        38007 => X"B8",  -- 184
        38008 => X"C3",  -- 195
        38009 => X"C0",  -- 192
        38010 => X"B8",  -- 184
        38011 => X"BE",  -- 190
        38012 => X"B7",  -- 183
        38013 => X"BB",  -- 187
        38014 => X"B6",  -- 182
        38015 => X"BA",  -- 186
        38016 => X"B2",  -- 178
        38017 => X"A4",  -- 164
        38018 => X"9B",  -- 155
        38019 => X"A8",  -- 168
        38020 => X"A8",  -- 168
        38021 => X"A4",  -- 164
        38022 => X"9D",  -- 157
        38023 => X"A0",  -- 160
        38024 => X"9B",  -- 155
        38025 => X"A1",  -- 161
        38026 => X"A1",  -- 161
        38027 => X"A3",  -- 163
        38028 => X"97",  -- 151
        38029 => X"9A",  -- 154
        38030 => X"9B",  -- 155
        38031 => X"92",  -- 146
        38032 => X"98",  -- 152
        38033 => X"94",  -- 148
        38034 => X"99",  -- 153
        38035 => X"9E",  -- 158
        38036 => X"91",  -- 145
        38037 => X"A1",  -- 161
        38038 => X"9B",  -- 155
        38039 => X"A4",  -- 164
        38040 => X"A0",  -- 160
        38041 => X"A7",  -- 167
        38042 => X"A4",  -- 164
        38043 => X"99",  -- 153
        38044 => X"9E",  -- 158
        38045 => X"AD",  -- 173
        38046 => X"B0",  -- 176
        38047 => X"A3",  -- 163
        38048 => X"AC",  -- 172
        38049 => X"B1",  -- 177
        38050 => X"AF",  -- 175
        38051 => X"B2",  -- 178
        38052 => X"C3",  -- 195
        38053 => X"C4",  -- 196
        38054 => X"BC",  -- 188
        38055 => X"C1",  -- 193
        38056 => X"B2",  -- 178
        38057 => X"9D",  -- 157
        38058 => X"94",  -- 148
        38059 => X"8C",  -- 140
        38060 => X"90",  -- 144
        38061 => X"91",  -- 145
        38062 => X"88",  -- 136
        38063 => X"98",  -- 152
        38064 => X"B8",  -- 184
        38065 => X"BE",  -- 190
        38066 => X"C2",  -- 194
        38067 => X"C0",  -- 192
        38068 => X"BB",  -- 187
        38069 => X"B7",  -- 183
        38070 => X"B4",  -- 180
        38071 => X"B2",  -- 178
        38072 => X"BD",  -- 189
        38073 => X"BD",  -- 189
        38074 => X"C0",  -- 192
        38075 => X"A9",  -- 169
        38076 => X"7A",  -- 122
        38077 => X"63",  -- 99
        38078 => X"66",  -- 102
        38079 => X"67",  -- 103
        38080 => X"45",  -- 69
        38081 => X"47",  -- 71
        38082 => X"4A",  -- 74
        38083 => X"4C",  -- 76
        38084 => X"4D",  -- 77
        38085 => X"4E",  -- 78
        38086 => X"4F",  -- 79
        38087 => X"50",  -- 80
        38088 => X"4E",  -- 78
        38089 => X"53",  -- 83
        38090 => X"57",  -- 87
        38091 => X"58",  -- 88
        38092 => X"54",  -- 84
        38093 => X"50",  -- 80
        38094 => X"4E",  -- 78
        38095 => X"4D",  -- 77
        38096 => X"47",  -- 71
        38097 => X"47",  -- 71
        38098 => X"49",  -- 73
        38099 => X"4D",  -- 77
        38100 => X"53",  -- 83
        38101 => X"55",  -- 85
        38102 => X"53",  -- 83
        38103 => X"51",  -- 81
        38104 => X"4C",  -- 76
        38105 => X"49",  -- 73
        38106 => X"55",  -- 85
        38107 => X"67",  -- 103
        38108 => X"6F",  -- 111
        38109 => X"79",  -- 121
        38110 => X"83",  -- 131
        38111 => X"89",  -- 137
        38112 => X"7D",  -- 125
        38113 => X"65",  -- 101
        38114 => X"48",  -- 72
        38115 => X"25",  -- 37
        38116 => X"14",  -- 20
        38117 => X"0F",  -- 15
        38118 => X"25",  -- 37
        38119 => X"63",  -- 99
        38120 => X"87",  -- 135
        38121 => X"93",  -- 147
        38122 => X"68",  -- 104
        38123 => X"1D",  -- 29
        38124 => X"0E",  -- 14
        38125 => X"29",  -- 41
        38126 => X"67",  -- 103
        38127 => X"7B",  -- 123
        38128 => X"71",  -- 113
        38129 => X"66",  -- 102
        38130 => X"24",  -- 36
        38131 => X"0B",  -- 11
        38132 => X"27",  -- 39
        38133 => X"47",  -- 71
        38134 => X"5D",  -- 93
        38135 => X"53",  -- 83
        38136 => X"38",  -- 56
        38137 => X"12",  -- 18
        38138 => X"18",  -- 24
        38139 => X"5C",  -- 92
        38140 => X"9A",  -- 154
        38141 => X"A5",  -- 165
        38142 => X"91",  -- 145
        38143 => X"7C",  -- 124
        38144 => X"45",  -- 69
        38145 => X"2B",  -- 43
        38146 => X"15",  -- 21
        38147 => X"12",  -- 18
        38148 => X"14",  -- 20
        38149 => X"13",  -- 19
        38150 => X"10",  -- 16
        38151 => X"11",  -- 17
        38152 => X"13",  -- 19
        38153 => X"0F",  -- 15
        38154 => X"02",  -- 2
        38155 => X"26",  -- 38
        38156 => X"85",  -- 133
        38157 => X"7C",  -- 124
        38158 => X"46",  -- 70
        38159 => X"35",  -- 53
        38160 => X"25",  -- 37
        38161 => X"29",  -- 41
        38162 => X"28",  -- 40
        38163 => X"27",  -- 39
        38164 => X"2F",  -- 47
        38165 => X"33",  -- 51
        38166 => X"37",  -- 55
        38167 => X"3F",  -- 63
        38168 => X"46",  -- 70
        38169 => X"4A",  -- 74
        38170 => X"4D",  -- 77
        38171 => X"4A",  -- 74
        38172 => X"4C",  -- 76
        38173 => X"3A",  -- 58
        38174 => X"5A",  -- 90
        38175 => X"51",  -- 81
        38176 => X"41",  -- 65
        38177 => X"45",  -- 69
        38178 => X"55",  -- 85
        38179 => X"54",  -- 84
        38180 => X"60",  -- 96
        38181 => X"4B",  -- 75
        38182 => X"4D",  -- 77
        38183 => X"51",  -- 81
        38184 => X"52",  -- 82
        38185 => X"49",  -- 73
        38186 => X"4B",  -- 75
        38187 => X"50",  -- 80
        38188 => X"43",  -- 67
        38189 => X"66",  -- 102
        38190 => X"89",  -- 137
        38191 => X"BB",  -- 187
        38192 => X"CE",  -- 206
        38193 => X"7B",  -- 123
        38194 => X"0B",  -- 11
        38195 => X"30",  -- 48
        38196 => X"27",  -- 39
        38197 => X"31",  -- 49
        38198 => X"1E",  -- 30
        38199 => X"21",  -- 33
        38200 => X"20",  -- 32
        38201 => X"17",  -- 23
        38202 => X"1C",  -- 28
        38203 => X"1E",  -- 30
        38204 => X"45",  -- 69
        38205 => X"82",  -- 130
        38206 => X"9A",  -- 154
        38207 => X"AD",  -- 173
        38208 => X"C0",  -- 192
        38209 => X"C0",  -- 192
        38210 => X"55",  -- 85
        38211 => X"11",  -- 17
        38212 => X"2B",  -- 43
        38213 => X"41",  -- 65
        38214 => X"55",  -- 85
        38215 => X"6B",  -- 107
        38216 => X"75",  -- 117
        38217 => X"7B",  -- 123
        38218 => X"A4",  -- 164
        38219 => X"B6",  -- 182
        38220 => X"B7",  -- 183
        38221 => X"B8",  -- 184
        38222 => X"AF",  -- 175
        38223 => X"C0",  -- 192
        38224 => X"B7",  -- 183
        38225 => X"A3",  -- 163
        38226 => X"2E",  -- 46
        38227 => X"16",  -- 22
        38228 => X"3B",  -- 59
        38229 => X"B8",  -- 184
        38230 => X"D4",  -- 212
        38231 => X"CF",  -- 207
        38232 => X"CD",  -- 205
        38233 => X"D7",  -- 215
        38234 => X"9F",  -- 159
        38235 => X"25",  -- 37
        38236 => X"0D",  -- 13
        38237 => X"2A",  -- 42
        38238 => X"5D",  -- 93
        38239 => X"83",  -- 131
        38240 => X"A6",  -- 166
        38241 => X"A9",  -- 169
        38242 => X"B4",  -- 180
        38243 => X"C1",  -- 193
        38244 => X"C1",  -- 193
        38245 => X"B6",  -- 182
        38246 => X"B0",  -- 176
        38247 => X"B4",  -- 180
        38248 => X"BA",  -- 186
        38249 => X"BF",  -- 191
        38250 => X"C8",  -- 200
        38251 => X"D1",  -- 209
        38252 => X"CF",  -- 207
        38253 => X"B8",  -- 184
        38254 => X"96",  -- 150
        38255 => X"7C",  -- 124
        38256 => X"77",  -- 119
        38257 => X"62",  -- 98
        38258 => X"4D",  -- 77
        38259 => X"48",  -- 72
        38260 => X"4E",  -- 78
        38261 => X"56",  -- 86
        38262 => X"5F",  -- 95
        38263 => X"64",  -- 100
        38264 => X"5E",  -- 94
        38265 => X"44",  -- 68
        38266 => X"3A",  -- 58
        38267 => X"45",  -- 69
        38268 => X"4C",  -- 76
        38269 => X"40",  -- 64
        38270 => X"34",  -- 52
        38271 => X"35",  -- 53
        38272 => X"31",  -- 49
        38273 => X"3A",  -- 58
        38274 => X"41",  -- 65
        38275 => X"47",  -- 71
        38276 => X"54",  -- 84
        38277 => X"65",  -- 101
        38278 => X"6A",  -- 106
        38279 => X"66",  -- 102
        38280 => X"79",  -- 121
        38281 => X"82",  -- 130
        38282 => X"83",  -- 131
        38283 => X"83",  -- 131
        38284 => X"84",  -- 132
        38285 => X"7B",  -- 123
        38286 => X"78",  -- 120
        38287 => X"7E",  -- 126
        38288 => X"81",  -- 129
        38289 => X"7D",  -- 125
        38290 => X"85",  -- 133
        38291 => X"90",  -- 144
        38292 => X"8B",  -- 139
        38293 => X"79",  -- 121
        38294 => X"77",  -- 119
        38295 => X"83",  -- 131
        38296 => X"84",  -- 132
        38297 => X"77",  -- 119
        38298 => X"6D",  -- 109
        38299 => X"6D",  -- 109
        38300 => X"6B",  -- 107
        38301 => X"64",  -- 100
        38302 => X"60",  -- 96
        38303 => X"63",  -- 99
        38304 => X"5F",  -- 95
        38305 => X"5C",  -- 92
        38306 => X"5D",  -- 93
        38307 => X"61",  -- 97
        38308 => X"5E",  -- 94
        38309 => X"55",  -- 85
        38310 => X"4E",  -- 78
        38311 => X"4C",  -- 76
        38312 => X"49",  -- 73
        38313 => X"42",  -- 66
        38314 => X"40",  -- 64
        38315 => X"49",  -- 73
        38316 => X"50",  -- 80
        38317 => X"50",  -- 80
        38318 => X"4C",  -- 76
        38319 => X"4A",  -- 74
        38320 => X"63",  -- 99
        38321 => X"88",  -- 136
        38322 => X"9E",  -- 158
        38323 => X"AC",  -- 172
        38324 => X"AC",  -- 172
        38325 => X"AD",  -- 173
        38326 => X"BC",  -- 188
        38327 => X"BB",  -- 187
        38328 => X"BE",  -- 190
        38329 => X"B7",  -- 183
        38330 => X"B5",  -- 181
        38331 => X"BE",  -- 190
        38332 => X"C1",  -- 193
        38333 => X"BD",  -- 189
        38334 => X"B5",  -- 181
        38335 => X"B4",  -- 180
        38336 => X"B7",  -- 183
        38337 => X"AC",  -- 172
        38338 => X"9D",  -- 157
        38339 => X"AB",  -- 171
        38340 => X"A5",  -- 165
        38341 => X"A9",  -- 169
        38342 => X"A1",  -- 161
        38343 => X"AB",  -- 171
        38344 => X"9C",  -- 156
        38345 => X"A6",  -- 166
        38346 => X"9E",  -- 158
        38347 => X"A6",  -- 166
        38348 => X"94",  -- 148
        38349 => X"9E",  -- 158
        38350 => X"9A",  -- 154
        38351 => X"8F",  -- 143
        38352 => X"9B",  -- 155
        38353 => X"95",  -- 149
        38354 => X"9B",  -- 155
        38355 => X"A2",  -- 162
        38356 => X"97",  -- 151
        38357 => X"A5",  -- 165
        38358 => X"9F",  -- 159
        38359 => X"A8",  -- 168
        38360 => X"A7",  -- 167
        38361 => X"9E",  -- 158
        38362 => X"9A",  -- 154
        38363 => X"A3",  -- 163
        38364 => X"A8",  -- 168
        38365 => X"A8",  -- 168
        38366 => X"AC",  -- 172
        38367 => X"B6",  -- 182
        38368 => X"B7",  -- 183
        38369 => X"BB",  -- 187
        38370 => X"B2",  -- 178
        38371 => X"B8",  -- 184
        38372 => X"CB",  -- 203
        38373 => X"CD",  -- 205
        38374 => X"C1",  -- 193
        38375 => X"C4",  -- 196
        38376 => X"C2",  -- 194
        38377 => X"A8",  -- 168
        38378 => X"91",  -- 145
        38379 => X"7A",  -- 122
        38380 => X"8D",  -- 141
        38381 => X"A0",  -- 160
        38382 => X"9B",  -- 155
        38383 => X"AD",  -- 173
        38384 => X"AC",  -- 172
        38385 => X"BC",  -- 188
        38386 => X"C4",  -- 196
        38387 => X"B9",  -- 185
        38388 => X"AB",  -- 171
        38389 => X"A8",  -- 168
        38390 => X"AC",  -- 172
        38391 => X"AE",  -- 174
        38392 => X"BB",  -- 187
        38393 => X"B6",  -- 182
        38394 => X"BD",  -- 189
        38395 => X"AC",  -- 172
        38396 => X"74",  -- 116
        38397 => X"4F",  -- 79
        38398 => X"56",  -- 86
        38399 => X"64",  -- 100
        38400 => X"44",  -- 68
        38401 => X"42",  -- 66
        38402 => X"40",  -- 64
        38403 => X"42",  -- 66
        38404 => X"47",  -- 71
        38405 => X"4B",  -- 75
        38406 => X"4D",  -- 77
        38407 => X"4D",  -- 77
        38408 => X"4D",  -- 77
        38409 => X"4E",  -- 78
        38410 => X"50",  -- 80
        38411 => X"52",  -- 82
        38412 => X"53",  -- 83
        38413 => X"51",  -- 81
        38414 => X"4E",  -- 78
        38415 => X"4A",  -- 74
        38416 => X"47",  -- 71
        38417 => X"49",  -- 73
        38418 => X"4C",  -- 76
        38419 => X"50",  -- 80
        38420 => X"54",  -- 84
        38421 => X"56",  -- 86
        38422 => X"53",  -- 83
        38423 => X"53",  -- 83
        38424 => X"55",  -- 85
        38425 => X"49",  -- 73
        38426 => X"50",  -- 80
        38427 => X"72",  -- 114
        38428 => X"70",  -- 112
        38429 => X"72",  -- 114
        38430 => X"92",  -- 146
        38431 => X"83",  -- 131
        38432 => X"87",  -- 135
        38433 => X"67",  -- 103
        38434 => X"4E",  -- 78
        38435 => X"27",  -- 39
        38436 => X"18",  -- 24
        38437 => X"12",  -- 18
        38438 => X"1D",  -- 29
        38439 => X"6E",  -- 110
        38440 => X"89",  -- 137
        38441 => X"9A",  -- 154
        38442 => X"71",  -- 113
        38443 => X"1B",  -- 27
        38444 => X"13",  -- 19
        38445 => X"19",  -- 25
        38446 => X"64",  -- 100
        38447 => X"7A",  -- 122
        38448 => X"6F",  -- 111
        38449 => X"3E",  -- 62
        38450 => X"2D",  -- 45
        38451 => X"19",  -- 25
        38452 => X"3A",  -- 58
        38453 => X"4E",  -- 78
        38454 => X"51",  -- 81
        38455 => X"54",  -- 84
        38456 => X"4D",  -- 77
        38457 => X"4D",  -- 77
        38458 => X"34",  -- 52
        38459 => X"1E",  -- 30
        38460 => X"48",  -- 72
        38461 => X"93",  -- 147
        38462 => X"AE",  -- 174
        38463 => X"95",  -- 149
        38464 => X"7C",  -- 124
        38465 => X"5B",  -- 91
        38466 => X"3D",  -- 61
        38467 => X"24",  -- 36
        38468 => X"1A",  -- 26
        38469 => X"17",  -- 23
        38470 => X"0C",  -- 12
        38471 => X"09",  -- 9
        38472 => X"12",  -- 18
        38473 => X"06",  -- 6
        38474 => X"0E",  -- 14
        38475 => X"0B",  -- 11
        38476 => X"62",  -- 98
        38477 => X"7A",  -- 122
        38478 => X"42",  -- 66
        38479 => X"3A",  -- 58
        38480 => X"2B",  -- 43
        38481 => X"2A",  -- 42
        38482 => X"29",  -- 41
        38483 => X"28",  -- 40
        38484 => X"2A",  -- 42
        38485 => X"31",  -- 49
        38486 => X"36",  -- 54
        38487 => X"3C",  -- 60
        38488 => X"4B",  -- 75
        38489 => X"47",  -- 71
        38490 => X"56",  -- 86
        38491 => X"4B",  -- 75
        38492 => X"47",  -- 71
        38493 => X"3A",  -- 58
        38494 => X"4C",  -- 76
        38495 => X"51",  -- 81
        38496 => X"4D",  -- 77
        38497 => X"5D",  -- 93
        38498 => X"52",  -- 82
        38499 => X"4F",  -- 79
        38500 => X"53",  -- 83
        38501 => X"51",  -- 81
        38502 => X"4E",  -- 78
        38503 => X"41",  -- 65
        38504 => X"43",  -- 67
        38505 => X"45",  -- 69
        38506 => X"56",  -- 86
        38507 => X"49",  -- 73
        38508 => X"45",  -- 69
        38509 => X"61",  -- 97
        38510 => X"7C",  -- 124
        38511 => X"A5",  -- 165
        38512 => X"AF",  -- 175
        38513 => X"4D",  -- 77
        38514 => X"10",  -- 16
        38515 => X"20",  -- 32
        38516 => X"3B",  -- 59
        38517 => X"2B",  -- 43
        38518 => X"0A",  -- 10
        38519 => X"27",  -- 39
        38520 => X"26",  -- 38
        38521 => X"1F",  -- 31
        38522 => X"3B",  -- 59
        38523 => X"4F",  -- 79
        38524 => X"78",  -- 120
        38525 => X"AF",  -- 175
        38526 => X"B7",  -- 183
        38527 => X"BC",  -- 188
        38528 => X"A1",  -- 161
        38529 => X"3F",  -- 63
        38530 => X"0A",  -- 10
        38531 => X"2C",  -- 44
        38532 => X"51",  -- 81
        38533 => X"56",  -- 86
        38534 => X"66",  -- 102
        38535 => X"83",  -- 131
        38536 => X"83",  -- 131
        38537 => X"90",  -- 144
        38538 => X"9B",  -- 155
        38539 => X"A6",  -- 166
        38540 => X"AE",  -- 174
        38541 => X"7D",  -- 125
        38542 => X"B0",  -- 176
        38543 => X"CA",  -- 202
        38544 => X"B8",  -- 184
        38545 => X"9C",  -- 156
        38546 => X"38",  -- 56
        38547 => X"13",  -- 19
        38548 => X"4B",  -- 75
        38549 => X"C5",  -- 197
        38550 => X"D2",  -- 210
        38551 => X"CF",  -- 207
        38552 => X"CD",  -- 205
        38553 => X"D2",  -- 210
        38554 => X"A1",  -- 161
        38555 => X"2C",  -- 44
        38556 => X"10",  -- 16
        38557 => X"28",  -- 40
        38558 => X"61",  -- 97
        38559 => X"95",  -- 149
        38560 => X"A3",  -- 163
        38561 => X"AE",  -- 174
        38562 => X"BF",  -- 191
        38563 => X"C7",  -- 199
        38564 => X"AA",  -- 170
        38565 => X"AC",  -- 172
        38566 => X"A4",  -- 164
        38567 => X"B1",  -- 177
        38568 => X"C0",  -- 192
        38569 => X"BA",  -- 186
        38570 => X"C9",  -- 201
        38571 => X"CE",  -- 206
        38572 => X"C2",  -- 194
        38573 => X"BE",  -- 190
        38574 => X"A6",  -- 166
        38575 => X"74",  -- 116
        38576 => X"57",  -- 87
        38577 => X"5A",  -- 90
        38578 => X"55",  -- 85
        38579 => X"4B",  -- 75
        38580 => X"4E",  -- 78
        38581 => X"5D",  -- 93
        38582 => X"65",  -- 101
        38583 => X"62",  -- 98
        38584 => X"6B",  -- 107
        38585 => X"5F",  -- 95
        38586 => X"40",  -- 64
        38587 => X"22",  -- 34
        38588 => X"2B",  -- 43
        38589 => X"45",  -- 69
        38590 => X"40",  -- 64
        38591 => X"26",  -- 38
        38592 => X"25",  -- 37
        38593 => X"34",  -- 52
        38594 => X"40",  -- 64
        38595 => X"4A",  -- 74
        38596 => X"5D",  -- 93
        38597 => X"71",  -- 113
        38598 => X"6B",  -- 107
        38599 => X"58",  -- 88
        38600 => X"6F",  -- 111
        38601 => X"78",  -- 120
        38602 => X"80",  -- 128
        38603 => X"83",  -- 131
        38604 => X"7F",  -- 127
        38605 => X"7A",  -- 122
        38606 => X"78",  -- 120
        38607 => X"7A",  -- 122
        38608 => X"7D",  -- 125
        38609 => X"79",  -- 121
        38610 => X"79",  -- 121
        38611 => X"7F",  -- 127
        38612 => X"86",  -- 134
        38613 => X"84",  -- 132
        38614 => X"78",  -- 120
        38615 => X"6D",  -- 109
        38616 => X"78",  -- 120
        38617 => X"75",  -- 117
        38618 => X"6B",  -- 107
        38619 => X"63",  -- 99
        38620 => X"61",  -- 97
        38621 => X"64",  -- 100
        38622 => X"61",  -- 97
        38623 => X"5C",  -- 92
        38624 => X"5A",  -- 90
        38625 => X"58",  -- 88
        38626 => X"55",  -- 85
        38627 => X"54",  -- 84
        38628 => X"57",  -- 87
        38629 => X"59",  -- 89
        38630 => X"52",  -- 82
        38631 => X"48",  -- 72
        38632 => X"46",  -- 70
        38633 => X"42",  -- 66
        38634 => X"45",  -- 69
        38635 => X"55",  -- 85
        38636 => X"66",  -- 102
        38637 => X"69",  -- 105
        38638 => X"5D",  -- 93
        38639 => X"50",  -- 80
        38640 => X"65",  -- 101
        38641 => X"88",  -- 136
        38642 => X"A6",  -- 166
        38643 => X"B2",  -- 178
        38644 => X"B9",  -- 185
        38645 => X"BB",  -- 187
        38646 => X"B9",  -- 185
        38647 => X"BD",  -- 189
        38648 => X"BC",  -- 188
        38649 => X"B1",  -- 177
        38650 => X"AC",  -- 172
        38651 => X"BB",  -- 187
        38652 => X"C7",  -- 199
        38653 => X"BC",  -- 188
        38654 => X"B2",  -- 178
        38655 => X"BA",  -- 186
        38656 => X"B8",  -- 184
        38657 => X"A9",  -- 169
        38658 => X"A0",  -- 160
        38659 => X"B5",  -- 181
        38660 => X"B8",  -- 184
        38661 => X"A7",  -- 167
        38662 => X"A7",  -- 167
        38663 => X"A9",  -- 169
        38664 => X"A6",  -- 166
        38665 => X"93",  -- 147
        38666 => X"A3",  -- 163
        38667 => X"A2",  -- 162
        38668 => X"93",  -- 147
        38669 => X"9B",  -- 155
        38670 => X"A0",  -- 160
        38671 => X"98",  -- 152
        38672 => X"9D",  -- 157
        38673 => X"91",  -- 145
        38674 => X"9D",  -- 157
        38675 => X"AC",  -- 172
        38676 => X"A3",  -- 163
        38677 => X"9C",  -- 156
        38678 => X"A3",  -- 163
        38679 => X"A5",  -- 165
        38680 => X"AA",  -- 170
        38681 => X"AD",  -- 173
        38682 => X"A4",  -- 164
        38683 => X"A1",  -- 161
        38684 => X"AB",  -- 171
        38685 => X"A9",  -- 169
        38686 => X"A7",  -- 167
        38687 => X"B6",  -- 182
        38688 => X"B6",  -- 182
        38689 => X"B7",  -- 183
        38690 => X"BA",  -- 186
        38691 => X"BE",  -- 190
        38692 => X"C5",  -- 197
        38693 => X"C8",  -- 200
        38694 => X"C7",  -- 199
        38695 => X"C5",  -- 197
        38696 => X"C2",  -- 194
        38697 => X"AD",  -- 173
        38698 => X"95",  -- 149
        38699 => X"84",  -- 132
        38700 => X"80",  -- 128
        38701 => X"88",  -- 136
        38702 => X"A2",  -- 162
        38703 => X"BA",  -- 186
        38704 => X"B4",  -- 180
        38705 => X"B5",  -- 181
        38706 => X"C0",  -- 192
        38707 => X"BF",  -- 191
        38708 => X"A7",  -- 167
        38709 => X"98",  -- 152
        38710 => X"A2",  -- 162
        38711 => X"AD",  -- 173
        38712 => X"B6",  -- 182
        38713 => X"BA",  -- 186
        38714 => X"B8",  -- 184
        38715 => X"A5",  -- 165
        38716 => X"80",  -- 128
        38717 => X"58",  -- 88
        38718 => X"49",  -- 73
        38719 => X"4F",  -- 79
        38720 => X"41",  -- 65
        38721 => X"3F",  -- 63
        38722 => X"3E",  -- 62
        38723 => X"3F",  -- 63
        38724 => X"43",  -- 67
        38725 => X"47",  -- 71
        38726 => X"49",  -- 73
        38727 => X"49",  -- 73
        38728 => X"50",  -- 80
        38729 => X"50",  -- 80
        38730 => X"4F",  -- 79
        38731 => X"4F",  -- 79
        38732 => X"4F",  -- 79
        38733 => X"4E",  -- 78
        38734 => X"4C",  -- 76
        38735 => X"4B",  -- 75
        38736 => X"4A",  -- 74
        38737 => X"4B",  -- 75
        38738 => X"4E",  -- 78
        38739 => X"50",  -- 80
        38740 => X"55",  -- 85
        38741 => X"55",  -- 85
        38742 => X"53",  -- 83
        38743 => X"52",  -- 82
        38744 => X"4B",  -- 75
        38745 => X"50",  -- 80
        38746 => X"5A",  -- 90
        38747 => X"5A",  -- 90
        38748 => X"65",  -- 101
        38749 => X"7B",  -- 123
        38750 => X"85",  -- 133
        38751 => X"82",  -- 130
        38752 => X"7F",  -- 127
        38753 => X"5E",  -- 94
        38754 => X"4A",  -- 74
        38755 => X"27",  -- 39
        38756 => X"18",  -- 24
        38757 => X"12",  -- 18
        38758 => X"24",  -- 36
        38759 => X"75",  -- 117
        38760 => X"88",  -- 136
        38761 => X"93",  -- 147
        38762 => X"6B",  -- 107
        38763 => X"18",  -- 24
        38764 => X"0D",  -- 13
        38765 => X"1A",  -- 26
        38766 => X"69",  -- 105
        38767 => X"75",  -- 117
        38768 => X"6F",  -- 111
        38769 => X"36",  -- 54
        38770 => X"24",  -- 36
        38771 => X"1F",  -- 31
        38772 => X"41",  -- 65
        38773 => X"4A",  -- 74
        38774 => X"45",  -- 69
        38775 => X"48",  -- 72
        38776 => X"3C",  -- 60
        38777 => X"41",  -- 65
        38778 => X"3F",  -- 63
        38779 => X"31",  -- 49
        38780 => X"2C",  -- 44
        38781 => X"47",  -- 71
        38782 => X"7B",  -- 123
        38783 => X"A1",  -- 161
        38784 => X"A7",  -- 167
        38785 => X"88",  -- 136
        38786 => X"68",  -- 104
        38787 => X"4A",  -- 74
        38788 => X"37",  -- 55
        38789 => X"2A",  -- 42
        38790 => X"1C",  -- 28
        38791 => X"14",  -- 20
        38792 => X"13",  -- 19
        38793 => X"0F",  -- 15
        38794 => X"0E",  -- 14
        38795 => X"08",  -- 8
        38796 => X"52",  -- 82
        38797 => X"66",  -- 102
        38798 => X"3A",  -- 58
        38799 => X"2F",  -- 47
        38800 => X"2F",  -- 47
        38801 => X"2D",  -- 45
        38802 => X"2B",  -- 43
        38803 => X"2B",  -- 43
        38804 => X"2E",  -- 46
        38805 => X"34",  -- 52
        38806 => X"3D",  -- 61
        38807 => X"42",  -- 66
        38808 => X"40",  -- 64
        38809 => X"4E",  -- 78
        38810 => X"5D",  -- 93
        38811 => X"55",  -- 85
        38812 => X"53",  -- 83
        38813 => X"54",  -- 84
        38814 => X"52",  -- 82
        38815 => X"40",  -- 64
        38816 => X"53",  -- 83
        38817 => X"62",  -- 98
        38818 => X"59",  -- 89
        38819 => X"51",  -- 81
        38820 => X"51",  -- 81
        38821 => X"4C",  -- 76
        38822 => X"4D",  -- 77
        38823 => X"47",  -- 71
        38824 => X"46",  -- 70
        38825 => X"49",  -- 73
        38826 => X"50",  -- 80
        38827 => X"48",  -- 72
        38828 => X"47",  -- 71
        38829 => X"59",  -- 89
        38830 => X"6F",  -- 111
        38831 => X"89",  -- 137
        38832 => X"85",  -- 133
        38833 => X"2C",  -- 44
        38834 => X"05",  -- 5
        38835 => X"1F",  -- 31
        38836 => X"26",  -- 38
        38837 => X"16",  -- 22
        38838 => X"1A",  -- 26
        38839 => X"34",  -- 52
        38840 => X"59",  -- 89
        38841 => X"72",  -- 114
        38842 => X"71",  -- 113
        38843 => X"84",  -- 132
        38844 => X"A1",  -- 161
        38845 => X"B6",  -- 182
        38846 => X"BF",  -- 191
        38847 => X"9F",  -- 159
        38848 => X"44",  -- 68
        38849 => X"23",  -- 35
        38850 => X"26",  -- 38
        38851 => X"4A",  -- 74
        38852 => X"57",  -- 87
        38853 => X"4C",  -- 76
        38854 => X"52",  -- 82
        38855 => X"64",  -- 100
        38856 => X"88",  -- 136
        38857 => X"94",  -- 148
        38858 => X"A9",  -- 169
        38859 => X"AE",  -- 174
        38860 => X"A7",  -- 167
        38861 => X"76",  -- 118
        38862 => X"AC",  -- 172
        38863 => X"C5",  -- 197
        38864 => X"BF",  -- 191
        38865 => X"A9",  -- 169
        38866 => X"41",  -- 65
        38867 => X"11",  -- 17
        38868 => X"46",  -- 70
        38869 => X"BF",  -- 191
        38870 => X"D5",  -- 213
        38871 => X"D8",  -- 216
        38872 => X"D2",  -- 210
        38873 => X"D1",  -- 209
        38874 => X"A5",  -- 165
        38875 => X"35",  -- 53
        38876 => X"0B",  -- 11
        38877 => X"1E",  -- 30
        38878 => X"63",  -- 99
        38879 => X"A0",  -- 160
        38880 => X"B0",  -- 176
        38881 => X"B5",  -- 181
        38882 => X"BA",  -- 186
        38883 => X"BE",  -- 190
        38884 => X"A9",  -- 169
        38885 => X"9D",  -- 157
        38886 => X"9E",  -- 158
        38887 => X"A5",  -- 165
        38888 => X"BD",  -- 189
        38889 => X"C0",  -- 192
        38890 => X"CD",  -- 205
        38891 => X"CF",  -- 207
        38892 => X"C3",  -- 195
        38893 => X"B8",  -- 184
        38894 => X"9D",  -- 157
        38895 => X"75",  -- 117
        38896 => X"58",  -- 88
        38897 => X"56",  -- 86
        38898 => X"4F",  -- 79
        38899 => X"4B",  -- 75
        38900 => X"53",  -- 83
        38901 => X"63",  -- 99
        38902 => X"6C",  -- 108
        38903 => X"6A",  -- 106
        38904 => X"64",  -- 100
        38905 => X"63",  -- 99
        38906 => X"54",  -- 84
        38907 => X"33",  -- 51
        38908 => X"1A",  -- 26
        38909 => X"17",  -- 23
        38910 => X"26",  -- 38
        38911 => X"36",  -- 54
        38912 => X"29",  -- 41
        38913 => X"34",  -- 52
        38914 => X"3F",  -- 63
        38915 => X"46",  -- 70
        38916 => X"55",  -- 85
        38917 => X"66",  -- 102
        38918 => X"65",  -- 101
        38919 => X"5B",  -- 91
        38920 => X"63",  -- 99
        38921 => X"6D",  -- 109
        38922 => X"7A",  -- 122
        38923 => X"80",  -- 128
        38924 => X"81",  -- 129
        38925 => X"7D",  -- 125
        38926 => X"79",  -- 121
        38927 => X"78",  -- 120
        38928 => X"7C",  -- 124
        38929 => X"79",  -- 121
        38930 => X"76",  -- 118
        38931 => X"76",  -- 118
        38932 => X"77",  -- 119
        38933 => X"77",  -- 119
        38934 => X"74",  -- 116
        38935 => X"70",  -- 112
        38936 => X"6C",  -- 108
        38937 => X"72",  -- 114
        38938 => X"71",  -- 113
        38939 => X"67",  -- 103
        38940 => X"5E",  -- 94
        38941 => X"5B",  -- 91
        38942 => X"5C",  -- 92
        38943 => X"5D",  -- 93
        38944 => X"57",  -- 87
        38945 => X"55",  -- 85
        38946 => X"52",  -- 82
        38947 => X"51",  -- 81
        38948 => X"54",  -- 84
        38949 => X"56",  -- 86
        38950 => X"50",  -- 80
        38951 => X"45",  -- 69
        38952 => X"45",  -- 69
        38953 => X"48",  -- 72
        38954 => X"50",  -- 80
        38955 => X"61",  -- 97
        38956 => X"71",  -- 113
        38957 => X"75",  -- 117
        38958 => X"6D",  -- 109
        38959 => X"63",  -- 99
        38960 => X"6D",  -- 109
        38961 => X"91",  -- 145
        38962 => X"AC",  -- 172
        38963 => X"B4",  -- 180
        38964 => X"BC",  -- 188
        38965 => X"C0",  -- 192
        38966 => X"BC",  -- 188
        38967 => X"B9",  -- 185
        38968 => X"C3",  -- 195
        38969 => X"BA",  -- 186
        38970 => X"B2",  -- 178
        38971 => X"BB",  -- 187
        38972 => X"C6",  -- 198
        38973 => X"BF",  -- 191
        38974 => X"B4",  -- 180
        38975 => X"B7",  -- 183
        38976 => X"B8",  -- 184
        38977 => X"AF",  -- 175
        38978 => X"A4",  -- 164
        38979 => X"B5",  -- 181
        38980 => X"BA",  -- 186
        38981 => X"AA",  -- 170
        38982 => X"AA",  -- 170
        38983 => X"A8",  -- 168
        38984 => X"A9",  -- 169
        38985 => X"98",  -- 152
        38986 => X"A6",  -- 166
        38987 => X"A6",  -- 166
        38988 => X"96",  -- 150
        38989 => X"9C",  -- 156
        38990 => X"A0",  -- 160
        38991 => X"9E",  -- 158
        38992 => X"9E",  -- 158
        38993 => X"96",  -- 150
        38994 => X"9B",  -- 155
        38995 => X"A4",  -- 164
        38996 => X"A3",  -- 163
        38997 => X"9F",  -- 159
        38998 => X"A0",  -- 160
        38999 => X"A0",  -- 160
        39000 => X"9E",  -- 158
        39001 => X"A9",  -- 169
        39002 => X"A9",  -- 169
        39003 => X"A3",  -- 163
        39004 => X"A5",  -- 165
        39005 => X"AA",  -- 170
        39006 => X"AE",  -- 174
        39007 => X"B4",  -- 180
        39008 => X"BB",  -- 187
        39009 => X"BB",  -- 187
        39010 => X"BE",  -- 190
        39011 => X"C2",  -- 194
        39012 => X"C5",  -- 197
        39013 => X"C6",  -- 198
        39014 => X"C6",  -- 198
        39015 => X"C5",  -- 197
        39016 => X"C3",  -- 195
        39017 => X"B7",  -- 183
        39018 => X"9E",  -- 158
        39019 => X"83",  -- 131
        39020 => X"7D",  -- 125
        39021 => X"8D",  -- 141
        39022 => X"A0",  -- 160
        39023 => X"AC",  -- 172
        39024 => X"C5",  -- 197
        39025 => X"BD",  -- 189
        39026 => X"B8",  -- 184
        39027 => X"B0",  -- 176
        39028 => X"A5",  -- 165
        39029 => X"A0",  -- 160
        39030 => X"A1",  -- 161
        39031 => X"A0",  -- 160
        39032 => X"B9",  -- 185
        39033 => X"BC",  -- 188
        39034 => X"AC",  -- 172
        39035 => X"9B",  -- 155
        39036 => X"87",  -- 135
        39037 => X"5D",  -- 93
        39038 => X"48",  -- 72
        39039 => X"5A",  -- 90
        39040 => X"3D",  -- 61
        39041 => X"3B",  -- 59
        39042 => X"3A",  -- 58
        39043 => X"3B",  -- 59
        39044 => X"3D",  -- 61
        39045 => X"40",  -- 64
        39046 => X"42",  -- 66
        39047 => X"43",  -- 67
        39048 => X"4B",  -- 75
        39049 => X"4A",  -- 74
        39050 => X"49",  -- 73
        39051 => X"48",  -- 72
        39052 => X"47",  -- 71
        39053 => X"48",  -- 72
        39054 => X"48",  -- 72
        39055 => X"4A",  -- 74
        39056 => X"4B",  -- 75
        39057 => X"4B",  -- 75
        39058 => X"4D",  -- 77
        39059 => X"4F",  -- 79
        39060 => X"52",  -- 82
        39061 => X"52",  -- 82
        39062 => X"50",  -- 80
        39063 => X"4E",  -- 78
        39064 => X"46",  -- 70
        39065 => X"4D",  -- 77
        39066 => X"5A",  -- 90
        39067 => X"4D",  -- 77
        39068 => X"62",  -- 98
        39069 => X"7F",  -- 127
        39070 => X"7A",  -- 122
        39071 => X"8E",  -- 142
        39072 => X"81",  -- 129
        39073 => X"60",  -- 96
        39074 => X"48",  -- 72
        39075 => X"29",  -- 41
        39076 => X"15",  -- 21
        39077 => X"0A",  -- 10
        39078 => X"20",  -- 32
        39079 => X"70",  -- 112
        39080 => X"88",  -- 136
        39081 => X"90",  -- 144
        39082 => X"6C",  -- 108
        39083 => X"23",  -- 35
        39084 => X"0B",  -- 11
        39085 => X"20",  -- 32
        39086 => X"70",  -- 112
        39087 => X"6F",  -- 111
        39088 => X"71",  -- 113
        39089 => X"32",  -- 50
        39090 => X"16",  -- 22
        39091 => X"20",  -- 32
        39092 => X"45",  -- 69
        39093 => X"4D",  -- 77
        39094 => X"49",  -- 73
        39095 => X"4D",  -- 77
        39096 => X"25",  -- 37
        39097 => X"2C",  -- 44
        39098 => X"44",  -- 68
        39099 => X"50",  -- 80
        39100 => X"33",  -- 51
        39101 => X"1B",  -- 27
        39102 => X"2C",  -- 44
        39103 => X"4D",  -- 77
        39104 => X"85",  -- 133
        39105 => X"9D",  -- 157
        39106 => X"A2",  -- 162
        39107 => X"8E",  -- 142
        39108 => X"86",  -- 134
        39109 => X"89",  -- 137
        39110 => X"61",  -- 97
        39111 => X"1D",  -- 29
        39112 => X"0C",  -- 12
        39113 => X"19",  -- 25
        39114 => X"0A",  -- 10
        39115 => X"05",  -- 5
        39116 => X"3E",  -- 62
        39117 => X"4D",  -- 77
        39118 => X"39",  -- 57
        39119 => X"2C",  -- 44
        39120 => X"29",  -- 41
        39121 => X"28",  -- 40
        39122 => X"27",  -- 39
        39123 => X"27",  -- 39
        39124 => X"29",  -- 41
        39125 => X"31",  -- 49
        39126 => X"3C",  -- 60
        39127 => X"43",  -- 67
        39128 => X"40",  -- 64
        39129 => X"50",  -- 80
        39130 => X"55",  -- 85
        39131 => X"56",  -- 86
        39132 => X"52",  -- 82
        39133 => X"5E",  -- 94
        39134 => X"5C",  -- 92
        39135 => X"57",  -- 87
        39136 => X"50",  -- 80
        39137 => X"60",  -- 96
        39138 => X"59",  -- 89
        39139 => X"52",  -- 82
        39140 => X"4D",  -- 77
        39141 => X"45",  -- 69
        39142 => X"4A",  -- 74
        39143 => X"4C",  -- 76
        39144 => X"44",  -- 68
        39145 => X"4A",  -- 74
        39146 => X"46",  -- 70
        39147 => X"4C",  -- 76
        39148 => X"52",  -- 82
        39149 => X"5B",  -- 91
        39150 => X"6F",  -- 111
        39151 => X"77",  -- 119
        39152 => X"77",  -- 119
        39153 => X"23",  -- 35
        39154 => X"04",  -- 4
        39155 => X"29",  -- 41
        39156 => X"24",  -- 36
        39157 => X"17",  -- 23
        39158 => X"5E",  -- 94
        39159 => X"8E",  -- 142
        39160 => X"B1",  -- 177
        39161 => X"C3",  -- 195
        39162 => X"A2",  -- 162
        39163 => X"9A",  -- 154
        39164 => X"AF",  -- 175
        39165 => X"A8",  -- 168
        39166 => X"7A",  -- 122
        39167 => X"31",  -- 49
        39168 => X"19",  -- 25
        39169 => X"2D",  -- 45
        39170 => X"56",  -- 86
        39171 => X"6E",  -- 110
        39172 => X"64",  -- 100
        39173 => X"55",  -- 85
        39174 => X"5A",  -- 90
        39175 => X"64",  -- 100
        39176 => X"8D",  -- 141
        39177 => X"93",  -- 147
        39178 => X"99",  -- 153
        39179 => X"80",  -- 128
        39180 => X"69",  -- 105
        39181 => X"62",  -- 98
        39182 => X"B2",  -- 178
        39183 => X"C6",  -- 198
        39184 => X"C4",  -- 196
        39185 => X"B8",  -- 184
        39186 => X"4E",  -- 78
        39187 => X"16",  -- 22
        39188 => X"48",  -- 72
        39189 => X"BC",  -- 188
        39190 => X"D8",  -- 216
        39191 => X"DD",  -- 221
        39192 => X"D3",  -- 211
        39193 => X"CD",  -- 205
        39194 => X"AF",  -- 175
        39195 => X"4F",  -- 79
        39196 => X"0F",  -- 15
        39197 => X"13",  -- 19
        39198 => X"54",  -- 84
        39199 => X"97",  -- 151
        39200 => X"BA",  -- 186
        39201 => X"C0",  -- 192
        39202 => X"BC",  -- 188
        39203 => X"BF",  -- 191
        39204 => X"B2",  -- 178
        39205 => X"91",  -- 145
        39206 => X"98",  -- 152
        39207 => X"93",  -- 147
        39208 => X"B5",  -- 181
        39209 => X"C4",  -- 196
        39210 => X"D1",  -- 209
        39211 => X"CF",  -- 207
        39212 => X"C5",  -- 197
        39213 => X"B7",  -- 183
        39214 => X"95",  -- 149
        39215 => X"72",  -- 114
        39216 => X"60",  -- 96
        39217 => X"5A",  -- 90
        39218 => X"54",  -- 84
        39219 => X"57",  -- 87
        39220 => X"61",  -- 97
        39221 => X"68",  -- 104
        39222 => X"68",  -- 104
        39223 => X"65",  -- 101
        39224 => X"50",  -- 80
        39225 => X"4B",  -- 75
        39226 => X"4E",  -- 78
        39227 => X"4A",  -- 74
        39228 => X"34",  -- 52
        39229 => X"19",  -- 25
        39230 => X"1A",  -- 26
        39231 => X"2D",  -- 45
        39232 => X"35",  -- 53
        39233 => X"3C",  -- 60
        39234 => X"43",  -- 67
        39235 => X"48",  -- 72
        39236 => X"4F",  -- 79
        39237 => X"57",  -- 87
        39238 => X"5A",  -- 90
        39239 => X"5B",  -- 91
        39240 => X"5C",  -- 92
        39241 => X"66",  -- 102
        39242 => X"73",  -- 115
        39243 => X"7D",  -- 125
        39244 => X"80",  -- 128
        39245 => X"7C",  -- 124
        39246 => X"77",  -- 119
        39247 => X"73",  -- 115
        39248 => X"7A",  -- 122
        39249 => X"7A",  -- 122
        39250 => X"79",  -- 121
        39251 => X"76",  -- 118
        39252 => X"72",  -- 114
        39253 => X"70",  -- 112
        39254 => X"71",  -- 113
        39255 => X"72",  -- 114
        39256 => X"64",  -- 100
        39257 => X"6B",  -- 107
        39258 => X"6E",  -- 110
        39259 => X"68",  -- 104
        39260 => X"5E",  -- 94
        39261 => X"59",  -- 89
        39262 => X"59",  -- 89
        39263 => X"59",  -- 89
        39264 => X"52",  -- 82
        39265 => X"51",  -- 81
        39266 => X"4D",  -- 77
        39267 => X"4C",  -- 76
        39268 => X"4F",  -- 79
        39269 => X"51",  -- 81
        39270 => X"4A",  -- 74
        39271 => X"41",  -- 65
        39272 => X"44",  -- 68
        39273 => X"4B",  -- 75
        39274 => X"59",  -- 89
        39275 => X"6A",  -- 106
        39276 => X"77",  -- 119
        39277 => X"7C",  -- 124
        39278 => X"79",  -- 121
        39279 => X"74",  -- 116
        39280 => X"79",  -- 121
        39281 => X"9C",  -- 156
        39282 => X"B0",  -- 176
        39283 => X"B3",  -- 179
        39284 => X"BD",  -- 189
        39285 => X"C5",  -- 197
        39286 => X"BF",  -- 191
        39287 => X"B8",  -- 184
        39288 => X"C7",  -- 199
        39289 => X"C0",  -- 192
        39290 => X"B7",  -- 183
        39291 => X"BA",  -- 186
        39292 => X"C3",  -- 195
        39293 => X"C0",  -- 192
        39294 => X"B2",  -- 178
        39295 => X"AF",  -- 175
        39296 => X"B9",  -- 185
        39297 => X"B5",  -- 181
        39298 => X"AC",  -- 172
        39299 => X"B7",  -- 183
        39300 => X"BA",  -- 186
        39301 => X"AF",  -- 175
        39302 => X"B0",  -- 176
        39303 => X"A8",  -- 168
        39304 => X"AE",  -- 174
        39305 => X"9B",  -- 155
        39306 => X"A8",  -- 168
        39307 => X"A9",  -- 169
        39308 => X"9B",  -- 155
        39309 => X"9B",  -- 155
        39310 => X"9E",  -- 158
        39311 => X"A4",  -- 164
        39312 => X"A0",  -- 160
        39313 => X"A1",  -- 161
        39314 => X"9C",  -- 156
        39315 => X"9C",  -- 156
        39316 => X"A5",  -- 165
        39317 => X"A7",  -- 167
        39318 => X"A2",  -- 162
        39319 => X"A1",  -- 161
        39320 => X"96",  -- 150
        39321 => X"A2",  -- 162
        39322 => X"AC",  -- 172
        39323 => X"A5",  -- 165
        39324 => X"A1",  -- 161
        39325 => X"AD",  -- 173
        39326 => X"B7",  -- 183
        39327 => X"B2",  -- 178
        39328 => X"BF",  -- 191
        39329 => X"C1",  -- 193
        39330 => X"C5",  -- 197
        39331 => X"C6",  -- 198
        39332 => X"C6",  -- 198
        39333 => X"C5",  -- 197
        39334 => X"C4",  -- 196
        39335 => X"C4",  -- 196
        39336 => X"C2",  -- 194
        39337 => X"C1",  -- 193
        39338 => X"AA",  -- 170
        39339 => X"86",  -- 134
        39340 => X"7E",  -- 126
        39341 => X"93",  -- 147
        39342 => X"A2",  -- 162
        39343 => X"A1",  -- 161
        39344 => X"BC",  -- 188
        39345 => X"C3",  -- 195
        39346 => X"C5",  -- 197
        39347 => X"B4",  -- 180
        39348 => X"9A",  -- 154
        39349 => X"8E",  -- 142
        39350 => X"94",  -- 148
        39351 => X"A0",  -- 160
        39352 => X"AF",  -- 175
        39353 => X"BD",  -- 189
        39354 => X"AB",  -- 171
        39355 => X"92",  -- 146
        39356 => X"85",  -- 133
        39357 => X"65",  -- 101
        39358 => X"4B",  -- 75
        39359 => X"54",  -- 84
        39360 => X"3E",  -- 62
        39361 => X"3C",  -- 60
        39362 => X"3A",  -- 58
        39363 => X"3A",  -- 58
        39364 => X"3A",  -- 58
        39365 => X"3C",  -- 60
        39366 => X"3D",  -- 61
        39367 => X"3E",  -- 62
        39368 => X"40",  -- 64
        39369 => X"41",  -- 65
        39370 => X"41",  -- 65
        39371 => X"41",  -- 65
        39372 => X"42",  -- 66
        39373 => X"43",  -- 67
        39374 => X"45",  -- 69
        39375 => X"46",  -- 70
        39376 => X"44",  -- 68
        39377 => X"45",  -- 69
        39378 => X"46",  -- 70
        39379 => X"48",  -- 72
        39380 => X"4A",  -- 74
        39381 => X"4B",  -- 75
        39382 => X"49",  -- 73
        39383 => X"48",  -- 72
        39384 => X"46",  -- 70
        39385 => X"41",  -- 65
        39386 => X"4E",  -- 78
        39387 => X"57",  -- 87
        39388 => X"67",  -- 103
        39389 => X"77",  -- 119
        39390 => X"80",  -- 128
        39391 => X"9C",  -- 156
        39392 => X"7F",  -- 127
        39393 => X"5D",  -- 93
        39394 => X"48",  -- 72
        39395 => X"2D",  -- 45
        39396 => X"13",  -- 19
        39397 => X"04",  -- 4
        39398 => X"1E",  -- 30
        39399 => X"68",  -- 104
        39400 => X"89",  -- 137
        39401 => X"91",  -- 145
        39402 => X"79",  -- 121
        39403 => X"38",  -- 56
        39404 => X"10",  -- 16
        39405 => X"28",  -- 40
        39406 => X"7C",  -- 124
        39407 => X"72",  -- 114
        39408 => X"78",  -- 120
        39409 => X"3A",  -- 58
        39410 => X"0E",  -- 14
        39411 => X"14",  -- 20
        39412 => X"3E",  -- 62
        39413 => X"58",  -- 88
        39414 => X"60",  -- 96
        39415 => X"65",  -- 101
        39416 => X"51",  -- 81
        39417 => X"46",  -- 70
        39418 => X"4D",  -- 77
        39419 => X"55",  -- 85
        39420 => X"46",  -- 70
        39421 => X"37",  -- 55
        39422 => X"33",  -- 51
        39423 => X"2F",  -- 47
        39424 => X"2E",  -- 46
        39425 => X"5A",  -- 90
        39426 => X"7E",  -- 126
        39427 => X"95",  -- 149
        39428 => X"B3",  -- 179
        39429 => X"C8",  -- 200
        39430 => X"94",  -- 148
        39431 => X"2D",  -- 45
        39432 => X"0D",  -- 13
        39433 => X"25",  -- 37
        39434 => X"0B",  -- 11
        39435 => X"06",  -- 6
        39436 => X"2B",  -- 43
        39437 => X"37",  -- 55
        39438 => X"35",  -- 53
        39439 => X"29",  -- 41
        39440 => X"22",  -- 34
        39441 => X"23",  -- 35
        39442 => X"24",  -- 36
        39443 => X"26",  -- 38
        39444 => X"29",  -- 41
        39445 => X"30",  -- 48
        39446 => X"38",  -- 56
        39447 => X"3F",  -- 63
        39448 => X"4A",  -- 74
        39449 => X"50",  -- 80
        39450 => X"4D",  -- 77
        39451 => X"59",  -- 89
        39452 => X"4F",  -- 79
        39453 => X"55",  -- 85
        39454 => X"56",  -- 86
        39455 => X"6F",  -- 111
        39456 => X"4E",  -- 78
        39457 => X"5F",  -- 95
        39458 => X"5A",  -- 90
        39459 => X"58",  -- 88
        39460 => X"54",  -- 84
        39461 => X"49",  -- 73
        39462 => X"4B",  -- 75
        39463 => X"4E",  -- 78
        39464 => X"49",  -- 73
        39465 => X"50",  -- 80
        39466 => X"44",  -- 68
        39467 => X"53",  -- 83
        39468 => X"5E",  -- 94
        39469 => X"61",  -- 97
        39470 => X"73",  -- 115
        39471 => X"6C",  -- 108
        39472 => X"63",  -- 99
        39473 => X"1E",  -- 30
        39474 => X"04",  -- 4
        39475 => X"2E",  -- 46
        39476 => X"2E",  -- 46
        39477 => X"15",  -- 21
        39478 => X"81",  -- 129
        39479 => X"D1",  -- 209
        39480 => X"DC",  -- 220
        39481 => X"D9",  -- 217
        39482 => X"B0",  -- 176
        39483 => X"5E",  -- 94
        39484 => X"47",  -- 71
        39485 => X"49",  -- 73
        39486 => X"25",  -- 37
        39487 => X"20",  -- 32
        39488 => X"3F",  -- 63
        39489 => X"4A",  -- 74
        39490 => X"58",  -- 88
        39491 => X"52",  -- 82
        39492 => X"40",  -- 64
        39493 => X"48",  -- 72
        39494 => X"6B",  -- 107
        39495 => X"86",  -- 134
        39496 => X"86",  -- 134
        39497 => X"7C",  -- 124
        39498 => X"6A",  -- 106
        39499 => X"33",  -- 51
        39500 => X"1F",  -- 31
        39501 => X"55",  -- 85
        39502 => X"B9",  -- 185
        39503 => X"BC",  -- 188
        39504 => X"C7",  -- 199
        39505 => X"C2",  -- 194
        39506 => X"58",  -- 88
        39507 => X"1F",  -- 31
        39508 => X"56",  -- 86
        39509 => X"BE",  -- 190
        39510 => X"DA",  -- 218
        39511 => X"D8",  -- 216
        39512 => X"D6",  -- 214
        39513 => X"CC",  -- 204
        39514 => X"BB",  -- 187
        39515 => X"70",  -- 112
        39516 => X"1F",  -- 31
        39517 => X"0F",  -- 15
        39518 => X"3F",  -- 63
        39519 => X"7E",  -- 126
        39520 => X"B7",  -- 183
        39521 => X"C8",  -- 200
        39522 => X"C5",  -- 197
        39523 => X"C9",  -- 201
        39524 => X"C2",  -- 194
        39525 => X"8D",  -- 141
        39526 => X"96",  -- 150
        39527 => X"8B",  -- 139
        39528 => X"A3",  -- 163
        39529 => X"C4",  -- 196
        39530 => X"D4",  -- 212
        39531 => X"CC",  -- 204
        39532 => X"C9",  -- 201
        39533 => X"BC",  -- 188
        39534 => X"91",  -- 145
        39535 => X"67",  -- 103
        39536 => X"5E",  -- 94
        39537 => X"5B",  -- 91
        39538 => X"5F",  -- 95
        39539 => X"69",  -- 105
        39540 => X"70",  -- 112
        39541 => X"6C",  -- 108
        39542 => X"64",  -- 100
        39543 => X"5E",  -- 94
        39544 => X"59",  -- 89
        39545 => X"3B",  -- 59
        39546 => X"2D",  -- 45
        39547 => X"34",  -- 52
        39548 => X"35",  -- 53
        39549 => X"27",  -- 39
        39550 => X"27",  -- 39
        39551 => X"36",  -- 54
        39552 => X"42",  -- 66
        39553 => X"47",  -- 71
        39554 => X"4E",  -- 78
        39555 => X"53",  -- 83
        39556 => X"51",  -- 81
        39557 => X"4F",  -- 79
        39558 => X"51",  -- 81
        39559 => X"57",  -- 87
        39560 => X"62",  -- 98
        39561 => X"66",  -- 102
        39562 => X"6F",  -- 111
        39563 => X"75",  -- 117
        39564 => X"78",  -- 120
        39565 => X"76",  -- 118
        39566 => X"71",  -- 113
        39567 => X"6E",  -- 110
        39568 => X"71",  -- 113
        39569 => X"75",  -- 117
        39570 => X"79",  -- 121
        39571 => X"79",  -- 121
        39572 => X"76",  -- 118
        39573 => X"71",  -- 113
        39574 => X"6D",  -- 109
        39575 => X"6C",  -- 108
        39576 => X"69",  -- 105
        39577 => X"67",  -- 103
        39578 => X"64",  -- 100
        39579 => X"63",  -- 99
        39580 => X"62",  -- 98
        39581 => X"5F",  -- 95
        39582 => X"59",  -- 89
        39583 => X"52",  -- 82
        39584 => X"4F",  -- 79
        39585 => X"4E",  -- 78
        39586 => X"4A",  -- 74
        39587 => X"48",  -- 72
        39588 => X"4B",  -- 75
        39589 => X"4C",  -- 76
        39590 => X"47",  -- 71
        39591 => X"40",  -- 64
        39592 => X"42",  -- 66
        39593 => X"51",  -- 81
        39594 => X"63",  -- 99
        39595 => X"71",  -- 113
        39596 => X"7A",  -- 122
        39597 => X"80",  -- 128
        39598 => X"83",  -- 131
        39599 => X"82",  -- 130
        39600 => X"86",  -- 134
        39601 => X"A5",  -- 165
        39602 => X"B3",  -- 179
        39603 => X"B0",  -- 176
        39604 => X"BB",  -- 187
        39605 => X"C6",  -- 198
        39606 => X"C2",  -- 194
        39607 => X"B9",  -- 185
        39608 => X"C0",  -- 192
        39609 => X"C1",  -- 193
        39610 => X"B9",  -- 185
        39611 => X"B6",  -- 182
        39612 => X"C0",  -- 192
        39613 => X"BE",  -- 190
        39614 => X"AF",  -- 175
        39615 => X"A8",  -- 168
        39616 => X"B5",  -- 181
        39617 => X"B7",  -- 183
        39618 => X"AE",  -- 174
        39619 => X"B6",  -- 182
        39620 => X"BB",  -- 187
        39621 => X"B4",  -- 180
        39622 => X"B5",  -- 181
        39623 => X"AD",  -- 173
        39624 => X"AF",  -- 175
        39625 => X"9D",  -- 157
        39626 => X"A8",  -- 168
        39627 => X"AA",  -- 170
        39628 => X"9E",  -- 158
        39629 => X"9A",  -- 154
        39630 => X"9B",  -- 155
        39631 => X"A8",  -- 168
        39632 => X"A4",  -- 164
        39633 => X"AD",  -- 173
        39634 => X"A3",  -- 163
        39635 => X"9D",  -- 157
        39636 => X"AB",  -- 171
        39637 => X"AF",  -- 175
        39638 => X"A8",  -- 168
        39639 => X"AA",  -- 170
        39640 => X"9A",  -- 154
        39641 => X"9C",  -- 156
        39642 => X"A7",  -- 167
        39643 => X"A8",  -- 168
        39644 => X"A1",  -- 161
        39645 => X"AF",  -- 175
        39646 => X"BC",  -- 188
        39647 => X"B5",  -- 181
        39648 => X"C2",  -- 194
        39649 => X"C5",  -- 197
        39650 => X"CA",  -- 202
        39651 => X"C9",  -- 201
        39652 => X"C6",  -- 198
        39653 => X"C4",  -- 196
        39654 => X"C2",  -- 194
        39655 => X"C2",  -- 194
        39656 => X"C1",  -- 193
        39657 => X"C2",  -- 194
        39658 => X"B0",  -- 176
        39659 => X"8F",  -- 143
        39660 => X"83",  -- 131
        39661 => X"91",  -- 145
        39662 => X"9F",  -- 159
        39663 => X"A1",  -- 161
        39664 => X"A7",  -- 167
        39665 => X"BE",  -- 190
        39666 => X"CD",  -- 205
        39667 => X"C0",  -- 192
        39668 => X"9B",  -- 155
        39669 => X"7B",  -- 123
        39670 => X"84",  -- 132
        39671 => X"A0",  -- 160
        39672 => X"A5",  -- 165
        39673 => X"BD",  -- 189
        39674 => X"BC",  -- 188
        39675 => X"9C",  -- 156
        39676 => X"80",  -- 128
        39677 => X"6B",  -- 107
        39678 => X"58",  -- 88
        39679 => X"4B",  -- 75
        39680 => X"41",  -- 65
        39681 => X"40",  -- 64
        39682 => X"3F",  -- 63
        39683 => X"3D",  -- 61
        39684 => X"3B",  -- 59
        39685 => X"3C",  -- 60
        39686 => X"3D",  -- 61
        39687 => X"3E",  -- 62
        39688 => X"3E",  -- 62
        39689 => X"40",  -- 64
        39690 => X"42",  -- 66
        39691 => X"42",  -- 66
        39692 => X"41",  -- 65
        39693 => X"40",  -- 64
        39694 => X"40",  -- 64
        39695 => X"41",  -- 65
        39696 => X"3E",  -- 62
        39697 => X"3E",  -- 62
        39698 => X"3E",  -- 62
        39699 => X"40",  -- 64
        39700 => X"42",  -- 66
        39701 => X"43",  -- 67
        39702 => X"42",  -- 66
        39703 => X"41",  -- 65
        39704 => X"42",  -- 66
        39705 => X"3C",  -- 60
        39706 => X"47",  -- 71
        39707 => X"64",  -- 100
        39708 => X"65",  -- 101
        39709 => X"6E",  -- 110
        39710 => X"90",  -- 144
        39711 => X"90",  -- 144
        39712 => X"6F",  -- 111
        39713 => X"54",  -- 84
        39714 => X"40",  -- 64
        39715 => X"2E",  -- 46
        39716 => X"14",  -- 20
        39717 => X"08",  -- 8
        39718 => X"27",  -- 39
        39719 => X"68",  -- 104
        39720 => X"86",  -- 134
        39721 => X"93",  -- 147
        39722 => X"82",  -- 130
        39723 => X"47",  -- 71
        39724 => X"12",  -- 18
        39725 => X"2A",  -- 42
        39726 => X"83",  -- 131
        39727 => X"84",  -- 132
        39728 => X"7C",  -- 124
        39729 => X"4A",  -- 74
        39730 => X"0F",  -- 15
        39731 => X"0A",  -- 10
        39732 => X"2C",  -- 44
        39733 => X"5A",  -- 90
        39734 => X"6D",  -- 109
        39735 => X"6B",  -- 107
        39736 => X"59",  -- 89
        39737 => X"42",  -- 66
        39738 => X"42",  -- 66
        39739 => X"4E",  -- 78
        39740 => X"4D",  -- 77
        39741 => X"51",  -- 81
        39742 => X"51",  -- 81
        39743 => X"42",  -- 66
        39744 => X"24",  -- 36
        39745 => X"1A",  -- 26
        39746 => X"2D",  -- 45
        39747 => X"73",  -- 115
        39748 => X"AE",  -- 174
        39749 => X"C1",  -- 193
        39750 => X"A1",  -- 161
        39751 => X"54",  -- 84
        39752 => X"14",  -- 20
        39753 => X"2F",  -- 47
        39754 => X"0E",  -- 14
        39755 => X"09",  -- 9
        39756 => X"1B",  -- 27
        39757 => X"21",  -- 33
        39758 => X"27",  -- 39
        39759 => X"1D",  -- 29
        39760 => X"20",  -- 32
        39761 => X"24",  -- 36
        39762 => X"28",  -- 40
        39763 => X"2B",  -- 43
        39764 => X"2F",  -- 47
        39765 => X"32",  -- 50
        39766 => X"39",  -- 57
        39767 => X"3E",  -- 62
        39768 => X"50",  -- 80
        39769 => X"57",  -- 87
        39770 => X"52",  -- 82
        39771 => X"61",  -- 97
        39772 => X"5A",  -- 90
        39773 => X"57",  -- 87
        39774 => X"48",  -- 72
        39775 => X"5B",  -- 91
        39776 => X"57",  -- 87
        39777 => X"63",  -- 99
        39778 => X"5F",  -- 95
        39779 => X"64",  -- 100
        39780 => X"64",  -- 100
        39781 => X"54",  -- 84
        39782 => X"50",  -- 80
        39783 => X"4E",  -- 78
        39784 => X"56",  -- 86
        39785 => X"58",  -- 88
        39786 => X"49",  -- 73
        39787 => X"54",  -- 84
        39788 => X"5D",  -- 93
        39789 => X"59",  -- 89
        39790 => X"61",  -- 97
        39791 => X"55",  -- 85
        39792 => X"41",  -- 65
        39793 => X"19",  -- 25
        39794 => X"04",  -- 4
        39795 => X"35",  -- 53
        39796 => X"46",  -- 70
        39797 => X"11",  -- 17
        39798 => X"74",  -- 116
        39799 => X"D4",  -- 212
        39800 => X"D9",  -- 217
        39801 => X"C7",  -- 199
        39802 => X"97",  -- 151
        39803 => X"46",  -- 70
        39804 => X"2D",  -- 45
        39805 => X"34",  -- 52
        39806 => X"2F",  -- 47
        39807 => X"50",  -- 80
        39808 => X"50",  -- 80
        39809 => X"41",  -- 65
        39810 => X"30",  -- 48
        39811 => X"1A",  -- 26
        39812 => X"0E",  -- 14
        39813 => X"23",  -- 35
        39814 => X"62",  -- 98
        39815 => X"93",  -- 147
        39816 => X"8E",  -- 142
        39817 => X"68",  -- 104
        39818 => X"48",  -- 72
        39819 => X"20",  -- 32
        39820 => X"1F",  -- 31
        39821 => X"6B",  -- 107
        39822 => X"C8",  -- 200
        39823 => X"C2",  -- 194
        39824 => X"CA",  -- 202
        39825 => X"C6",  -- 198
        39826 => X"56",  -- 86
        39827 => X"1D",  -- 29
        39828 => X"60",  -- 96
        39829 => X"C0",  -- 192
        39830 => X"DB",  -- 219
        39831 => X"D3",  -- 211
        39832 => X"DE",  -- 222
        39833 => X"CA",  -- 202
        39834 => X"B6",  -- 182
        39835 => X"7B",  -- 123
        39836 => X"2B",  -- 43
        39837 => X"14",  -- 20
        39838 => X"3A",  -- 58
        39839 => X"7B",  -- 123
        39840 => X"B0",  -- 176
        39841 => X"CE",  -- 206
        39842 => X"CD",  -- 205
        39843 => X"CE",  -- 206
        39844 => X"C8",  -- 200
        39845 => X"93",  -- 147
        39846 => X"9A",  -- 154
        39847 => X"8F",  -- 143
        39848 => X"93",  -- 147
        39849 => X"BF",  -- 191
        39850 => X"D2",  -- 210
        39851 => X"CA",  -- 202
        39852 => X"CB",  -- 203
        39853 => X"C4",  -- 196
        39854 => X"95",  -- 149
        39855 => X"60",  -- 96
        39856 => X"52",  -- 82
        39857 => X"56",  -- 86
        39858 => X"61",  -- 97
        39859 => X"6F",  -- 111
        39860 => X"75",  -- 117
        39861 => X"70",  -- 112
        39862 => X"69",  -- 105
        39863 => X"65",  -- 101
        39864 => X"59",  -- 89
        39865 => X"40",  -- 64
        39866 => X"2F",  -- 47
        39867 => X"2C",  -- 44
        39868 => X"2C",  -- 44
        39869 => X"27",  -- 39
        39870 => X"2B",  -- 43
        39871 => X"38",  -- 56
        39872 => X"45",  -- 69
        39873 => X"4B",  -- 75
        39874 => X"54",  -- 84
        39875 => X"5A",  -- 90
        39876 => X"58",  -- 88
        39877 => X"51",  -- 81
        39878 => X"50",  -- 80
        39879 => X"56",  -- 86
        39880 => X"69",  -- 105
        39881 => X"69",  -- 105
        39882 => X"6B",  -- 107
        39883 => X"6C",  -- 108
        39884 => X"6C",  -- 108
        39885 => X"6D",  -- 109
        39886 => X"6D",  -- 109
        39887 => X"6D",  -- 109
        39888 => X"6C",  -- 108
        39889 => X"6D",  -- 109
        39890 => X"70",  -- 112
        39891 => X"73",  -- 115
        39892 => X"73",  -- 115
        39893 => X"70",  -- 112
        39894 => X"69",  -- 105
        39895 => X"64",  -- 100
        39896 => X"6A",  -- 106
        39897 => X"65",  -- 101
        39898 => X"62",  -- 98
        39899 => X"61",  -- 97
        39900 => X"62",  -- 98
        39901 => X"5E",  -- 94
        39902 => X"59",  -- 89
        39903 => X"55",  -- 85
        39904 => X"4D",  -- 77
        39905 => X"4C",  -- 76
        39906 => X"49",  -- 73
        39907 => X"46",  -- 70
        39908 => X"47",  -- 71
        39909 => X"49",  -- 73
        39910 => X"47",  -- 71
        39911 => X"41",  -- 65
        39912 => X"44",  -- 68
        39913 => X"57",  -- 87
        39914 => X"6C",  -- 108
        39915 => X"78",  -- 120
        39916 => X"7D",  -- 125
        39917 => X"85",  -- 133
        39918 => X"8D",  -- 141
        39919 => X"92",  -- 146
        39920 => X"99",  -- 153
        39921 => X"B0",  -- 176
        39922 => X"B8",  -- 184
        39923 => X"B1",  -- 177
        39924 => X"BA",  -- 186
        39925 => X"C3",  -- 195
        39926 => X"C1",  -- 193
        39927 => X"BA",  -- 186
        39928 => X"BC",  -- 188
        39929 => X"BF",  -- 191
        39930 => X"BA",  -- 186
        39931 => X"B8",  -- 184
        39932 => X"C0",  -- 192
        39933 => X"C0",  -- 192
        39934 => X"B0",  -- 176
        39935 => X"A7",  -- 167
        39936 => X"AD",  -- 173
        39937 => X"B3",  -- 179
        39938 => X"AE",  -- 174
        39939 => X"B6",  -- 182
        39940 => X"BB",  -- 187
        39941 => X"B7",  -- 183
        39942 => X"BB",  -- 187
        39943 => X"B1",  -- 177
        39944 => X"B0",  -- 176
        39945 => X"A0",  -- 160
        39946 => X"A7",  -- 167
        39947 => X"AC",  -- 172
        39948 => X"A4",  -- 164
        39949 => X"9E",  -- 158
        39950 => X"9D",  -- 157
        39951 => X"AD",  -- 173
        39952 => X"A5",  -- 165
        39953 => X"B1",  -- 177
        39954 => X"A9",  -- 169
        39955 => X"A1",  -- 161
        39956 => X"AD",  -- 173
        39957 => X"B3",  -- 179
        39958 => X"B0",  -- 176
        39959 => X"B3",  -- 179
        39960 => X"AA",  -- 170
        39961 => X"9B",  -- 155
        39962 => X"A0",  -- 160
        39963 => X"A9",  -- 169
        39964 => X"A6",  -- 166
        39965 => X"AE",  -- 174
        39966 => X"BA",  -- 186
        39967 => X"BB",  -- 187
        39968 => X"C2",  -- 194
        39969 => X"C7",  -- 199
        39970 => X"CB",  -- 203
        39971 => X"CB",  -- 203
        39972 => X"C8",  -- 200
        39973 => X"C4",  -- 196
        39974 => X"C3",  -- 195
        39975 => X"C3",  -- 195
        39976 => X"BF",  -- 191
        39977 => X"BF",  -- 191
        39978 => X"B4",  -- 180
        39979 => X"9B",  -- 155
        39980 => X"89",  -- 137
        39981 => X"89",  -- 137
        39982 => X"96",  -- 150
        39983 => X"A0",  -- 160
        39984 => X"AD",  -- 173
        39985 => X"B1",  -- 177
        39986 => X"B5",  -- 181
        39987 => X"B8",  -- 184
        39988 => X"A8",  -- 168
        39989 => X"84",  -- 132
        39990 => X"7D",  -- 125
        39991 => X"94",  -- 148
        39992 => X"A9",  -- 169
        39993 => X"B1",  -- 177
        39994 => X"C1",  -- 193
        39995 => X"AF",  -- 175
        39996 => X"7E",  -- 126
        39997 => X"65",  -- 101
        39998 => X"63",  -- 99
        39999 => X"58",  -- 88
        40000 => X"46",  -- 70
        40001 => X"46",  -- 70
        40002 => X"45",  -- 69
        40003 => X"43",  -- 67
        40004 => X"41",  -- 65
        40005 => X"41",  -- 65
        40006 => X"44",  -- 68
        40007 => X"46",  -- 70
        40008 => X"48",  -- 72
        40009 => X"4A",  -- 74
        40010 => X"4B",  -- 75
        40011 => X"48",  -- 72
        40012 => X"43",  -- 67
        40013 => X"3F",  -- 63
        40014 => X"3E",  -- 62
        40015 => X"3F",  -- 63
        40016 => X"3C",  -- 60
        40017 => X"3C",  -- 60
        40018 => X"3B",  -- 59
        40019 => X"3C",  -- 60
        40020 => X"3E",  -- 62
        40021 => X"3E",  -- 62
        40022 => X"3D",  -- 61
        40023 => X"3D",  -- 61
        40024 => X"38",  -- 56
        40025 => X"41",  -- 65
        40026 => X"4C",  -- 76
        40027 => X"66",  -- 102
        40028 => X"5F",  -- 95
        40029 => X"6D",  -- 109
        40030 => X"92",  -- 146
        40031 => X"73",  -- 115
        40032 => X"68",  -- 104
        40033 => X"53",  -- 83
        40034 => X"40",  -- 64
        40035 => X"2F",  -- 47
        40036 => X"15",  -- 21
        40037 => X"0A",  -- 10
        40038 => X"29",  -- 41
        40039 => X"59",  -- 89
        40040 => X"82",  -- 130
        40041 => X"92",  -- 146
        40042 => X"84",  -- 132
        40043 => X"50",  -- 80
        40044 => X"13",  -- 19
        40045 => X"28",  -- 40
        40046 => X"82",  -- 130
        40047 => X"94",  -- 148
        40048 => X"77",  -- 119
        40049 => X"59",  -- 89
        40050 => X"18",  -- 24
        40051 => X"06",  -- 6
        40052 => X"1B",  -- 27
        40053 => X"4F",  -- 79
        40054 => X"67",  -- 103
        40055 => X"5E",  -- 94
        40056 => X"32",  -- 50
        40057 => X"11",  -- 17
        40058 => X"19",  -- 25
        40059 => X"3A",  -- 58
        40060 => X"42",  -- 66
        40061 => X"42",  -- 66
        40062 => X"3F",  -- 63
        40063 => X"2C",  -- 44
        40064 => X"37",  -- 55
        40065 => X"23",  -- 35
        40066 => X"26",  -- 38
        40067 => X"69",  -- 105
        40068 => X"A5",  -- 165
        40069 => X"C1",  -- 193
        40070 => X"B0",  -- 176
        40071 => X"60",  -- 96
        40072 => X"10",  -- 16
        40073 => X"24",  -- 36
        40074 => X"0A",  -- 10
        40075 => X"0C",  -- 12
        40076 => X"12",  -- 18
        40077 => X"19",  -- 25
        40078 => X"1E",  -- 30
        40079 => X"1C",  -- 28
        40080 => X"1E",  -- 30
        40081 => X"24",  -- 36
        40082 => X"2C",  -- 44
        40083 => X"2F",  -- 47
        40084 => X"32",  -- 50
        40085 => X"34",  -- 52
        40086 => X"38",  -- 56
        40087 => X"3C",  -- 60
        40088 => X"50",  -- 80
        40089 => X"5D",  -- 93
        40090 => X"52",  -- 82
        40091 => X"54",  -- 84
        40092 => X"61",  -- 97
        40093 => X"65",  -- 101
        40094 => X"50",  -- 80
        40095 => X"4E",  -- 78
        40096 => X"61",  -- 97
        40097 => X"67",  -- 103
        40098 => X"5F",  -- 95
        40099 => X"68",  -- 104
        40100 => X"6B",  -- 107
        40101 => X"5B",  -- 91
        40102 => X"52",  -- 82
        40103 => X"4F",  -- 79
        40104 => X"56",  -- 86
        40105 => X"55",  -- 85
        40106 => X"4E",  -- 78
        40107 => X"51",  -- 81
        40108 => X"53",  -- 83
        40109 => X"4D",  -- 77
        40110 => X"49",  -- 73
        40111 => X"40",  -- 64
        40112 => X"2F",  -- 47
        40113 => X"18",  -- 24
        40114 => X"05",  -- 5
        40115 => X"30",  -- 48
        40116 => X"4A",  -- 74
        40117 => X"1A",  -- 26
        40118 => X"77",  -- 119
        40119 => X"D2",  -- 210
        40120 => X"D1",  -- 209
        40121 => X"C0",  -- 192
        40122 => X"7E",  -- 126
        40123 => X"60",  -- 96
        40124 => X"5C",  -- 92
        40125 => X"4E",  -- 78
        40126 => X"56",  -- 86
        40127 => X"52",  -- 82
        40128 => X"32",  -- 50
        40129 => X"2E",  -- 46
        40130 => X"32",  -- 50
        40131 => X"31",  -- 49
        40132 => X"23",  -- 35
        40133 => X"2C",  -- 44
        40134 => X"5C",  -- 92
        40135 => X"87",  -- 135
        40136 => X"88",  -- 136
        40137 => X"3F",  -- 63
        40138 => X"16",  -- 22
        40139 => X"0E",  -- 14
        40140 => X"23",  -- 35
        40141 => X"70",  -- 112
        40142 => X"B8",  -- 184
        40143 => X"B8",  -- 184
        40144 => X"D0",  -- 208
        40145 => X"C7",  -- 199
        40146 => X"4D",  -- 77
        40147 => X"16",  -- 22
        40148 => X"68",  -- 104
        40149 => X"BF",  -- 191
        40150 => X"DD",  -- 221
        40151 => X"D3",  -- 211
        40152 => X"DE",  -- 222
        40153 => X"C4",  -- 196
        40154 => X"9F",  -- 159
        40155 => X"6B",  -- 107
        40156 => X"28",  -- 40
        40157 => X"15",  -- 21
        40158 => X"37",  -- 55
        40159 => X"80",  -- 128
        40160 => X"A8",  -- 168
        40161 => X"CE",  -- 206
        40162 => X"CE",  -- 206
        40163 => X"C9",  -- 201
        40164 => X"C2",  -- 194
        40165 => X"9D",  -- 157
        40166 => X"9C",  -- 156
        40167 => X"99",  -- 153
        40168 => X"92",  -- 146
        40169 => X"B4",  -- 180
        40170 => X"CC",  -- 204
        40171 => X"CD",  -- 205
        40172 => X"CB",  -- 203
        40173 => X"C5",  -- 197
        40174 => X"9C",  -- 156
        40175 => X"69",  -- 105
        40176 => X"59",  -- 89
        40177 => X"5E",  -- 94
        40178 => X"66",  -- 102
        40179 => X"6C",  -- 108
        40180 => X"6E",  -- 110
        40181 => X"6B",  -- 107
        40182 => X"67",  -- 103
        40183 => X"62",  -- 98
        40184 => X"57",  -- 87
        40185 => X"4B",  -- 75
        40186 => X"40",  -- 64
        40187 => X"3B",  -- 59
        40188 => X"3A",  -- 58
        40189 => X"38",  -- 56
        40190 => X"35",  -- 53
        40191 => X"34",  -- 52
        40192 => X"41",  -- 65
        40193 => X"49",  -- 73
        40194 => X"52",  -- 82
        40195 => X"5A",  -- 90
        40196 => X"5C",  -- 92
        40197 => X"59",  -- 89
        40198 => X"58",  -- 88
        40199 => X"5B",  -- 91
        40200 => X"6A",  -- 106
        40201 => X"69",  -- 105
        40202 => X"68",  -- 104
        40203 => X"66",  -- 102
        40204 => X"65",  -- 101
        40205 => X"67",  -- 103
        40206 => X"6C",  -- 108
        40207 => X"6F",  -- 111
        40208 => X"71",  -- 113
        40209 => X"6C",  -- 108
        40210 => X"68",  -- 104
        40211 => X"69",  -- 105
        40212 => X"6D",  -- 109
        40213 => X"6F",  -- 111
        40214 => X"6B",  -- 107
        40215 => X"66",  -- 102
        40216 => X"61",  -- 97
        40217 => X"63",  -- 99
        40218 => X"65",  -- 101
        40219 => X"62",  -- 98
        40220 => X"5A",  -- 90
        40221 => X"54",  -- 84
        40222 => X"55",  -- 85
        40223 => X"5B",  -- 91
        40224 => X"4E",  -- 78
        40225 => X"4C",  -- 76
        40226 => X"47",  -- 71
        40227 => X"43",  -- 67
        40228 => X"43",  -- 67
        40229 => X"47",  -- 71
        40230 => X"47",  -- 71
        40231 => X"43",  -- 67
        40232 => X"41",  -- 65
        40233 => X"57",  -- 87
        40234 => X"6D",  -- 109
        40235 => X"77",  -- 119
        40236 => X"7D",  -- 125
        40237 => X"89",  -- 137
        40238 => X"96",  -- 150
        40239 => X"9F",  -- 159
        40240 => X"A9",  -- 169
        40241 => X"BD",  -- 189
        40242 => X"C1",  -- 193
        40243 => X"B9",  -- 185
        40244 => X"BC",  -- 188
        40245 => X"C0",  -- 192
        40246 => X"BD",  -- 189
        40247 => X"BB",  -- 187
        40248 => X"BB",  -- 187
        40249 => X"C0",  -- 192
        40250 => X"BD",  -- 189
        40251 => X"BC",  -- 188
        40252 => X"C1",  -- 193
        40253 => X"BE",  -- 190
        40254 => X"B3",  -- 179
        40255 => X"B0",  -- 176
        40256 => X"A6",  -- 166
        40257 => X"AC",  -- 172
        40258 => X"A8",  -- 168
        40259 => X"B5",  -- 181
        40260 => X"BA",  -- 186
        40261 => X"B7",  -- 183
        40262 => X"BB",  -- 187
        40263 => X"B3",  -- 179
        40264 => X"AD",  -- 173
        40265 => X"A4",  -- 164
        40266 => X"A9",  -- 169
        40267 => X"AB",  -- 171
        40268 => X"AB",  -- 171
        40269 => X"A7",  -- 167
        40270 => X"A1",  -- 161
        40271 => X"AF",  -- 175
        40272 => X"A9",  -- 169
        40273 => X"AE",  -- 174
        40274 => X"AB",  -- 171
        40275 => X"A6",  -- 166
        40276 => X"AD",  -- 173
        40277 => X"B3",  -- 179
        40278 => X"B4",  -- 180
        40279 => X"B4",  -- 180
        40280 => X"B3",  -- 179
        40281 => X"A0",  -- 160
        40282 => X"9D",  -- 157
        40283 => X"A8",  -- 168
        40284 => X"AD",  -- 173
        40285 => X"AF",  -- 175
        40286 => X"B8",  -- 184
        40287 => X"C0",  -- 192
        40288 => X"C4",  -- 196
        40289 => X"C7",  -- 199
        40290 => X"CB",  -- 203
        40291 => X"CA",  -- 202
        40292 => X"C9",  -- 201
        40293 => X"C5",  -- 197
        40294 => X"C1",  -- 193
        40295 => X"BF",  -- 191
        40296 => X"BB",  -- 187
        40297 => X"B9",  -- 185
        40298 => X"B4",  -- 180
        40299 => X"A8",  -- 168
        40300 => X"94",  -- 148
        40301 => X"87",  -- 135
        40302 => X"8C",  -- 140
        40303 => X"99",  -- 153
        40304 => X"B0",  -- 176
        40305 => X"AC",  -- 172
        40306 => X"A4",  -- 164
        40307 => X"A6",  -- 166
        40308 => X"A3",  -- 163
        40309 => X"86",  -- 134
        40310 => X"79",  -- 121
        40311 => X"90",  -- 144
        40312 => X"AC",  -- 172
        40313 => X"9C",  -- 156
        40314 => X"AC",  -- 172
        40315 => X"AE",  -- 174
        40316 => X"7E",  -- 126
        40317 => X"56",  -- 86
        40318 => X"5C",  -- 92
        40319 => X"6A",  -- 106
        40320 => X"49",  -- 73
        40321 => X"4A",  -- 74
        40322 => X"4A",  -- 74
        40323 => X"49",  -- 73
        40324 => X"49",  -- 73
        40325 => X"4A",  -- 74
        40326 => X"4E",  -- 78
        40327 => X"51",  -- 81
        40328 => X"53",  -- 83
        40329 => X"54",  -- 84
        40330 => X"52",  -- 82
        40331 => X"4D",  -- 77
        40332 => X"46",  -- 70
        40333 => X"41",  -- 65
        40334 => X"41",  -- 65
        40335 => X"42",  -- 66
        40336 => X"42",  -- 66
        40337 => X"40",  -- 64
        40338 => X"3F",  -- 63
        40339 => X"3E",  -- 62
        40340 => X"3E",  -- 62
        40341 => X"3E",  -- 62
        40342 => X"3C",  -- 60
        40343 => X"3B",  -- 59
        40344 => X"36",  -- 54
        40345 => X"42",  -- 66
        40346 => X"53",  -- 83
        40347 => X"64",  -- 100
        40348 => X"67",  -- 103
        40349 => X"73",  -- 115
        40350 => X"7A",  -- 122
        40351 => X"66",  -- 102
        40352 => X"6D",  -- 109
        40353 => X"5A",  -- 90
        40354 => X"46",  -- 70
        40355 => X"32",  -- 50
        40356 => X"14",  -- 20
        40357 => X"08",  -- 8
        40358 => X"23",  -- 35
        40359 => X"40",  -- 64
        40360 => X"81",  -- 129
        40361 => X"97",  -- 151
        40362 => X"8C",  -- 140
        40363 => X"62",  -- 98
        40364 => X"21",  -- 33
        40365 => X"29",  -- 41
        40366 => X"77",  -- 119
        40367 => X"8E",  -- 142
        40368 => X"73",  -- 115
        40369 => X"61",  -- 97
        40370 => X"1E",  -- 30
        40371 => X"0A",  -- 10
        40372 => X"12",  -- 18
        40373 => X"47",  -- 71
        40374 => X"63",  -- 99
        40375 => X"5C",  -- 92
        40376 => X"44",  -- 68
        40377 => X"18",  -- 24
        40378 => X"15",  -- 21
        40379 => X"26",  -- 38
        40380 => X"23",  -- 35
        40381 => X"2D",  -- 45
        40382 => X"42",  -- 66
        40383 => X"3F",  -- 63
        40384 => X"3E",  -- 62
        40385 => X"44",  -- 68
        40386 => X"43",  -- 67
        40387 => X"64",  -- 100
        40388 => X"8B",  -- 139
        40389 => X"B3",  -- 179
        40390 => X"B0",  -- 176
        40391 => X"53",  -- 83
        40392 => X"07",  -- 7
        40393 => X"13",  -- 19
        40394 => X"04",  -- 4
        40395 => X"0E",  -- 14
        40396 => X"10",  -- 16
        40397 => X"1D",  -- 29
        40398 => X"1A",  -- 26
        40399 => X"20",  -- 32
        40400 => X"1E",  -- 30
        40401 => X"25",  -- 37
        40402 => X"2C",  -- 44
        40403 => X"2E",  -- 46
        40404 => X"2F",  -- 47
        40405 => X"30",  -- 48
        40406 => X"36",  -- 54
        40407 => X"3B",  -- 59
        40408 => X"4B",  -- 75
        40409 => X"58",  -- 88
        40410 => X"53",  -- 83
        40411 => X"4A",  -- 74
        40412 => X"60",  -- 96
        40413 => X"5E",  -- 94
        40414 => X"5A",  -- 90
        40415 => X"5E",  -- 94
        40416 => X"65",  -- 101
        40417 => X"66",  -- 102
        40418 => X"5C",  -- 92
        40419 => X"64",  -- 100
        40420 => X"69",  -- 105
        40421 => X"5C",  -- 92
        40422 => X"5A",  -- 90
        40423 => X"5B",  -- 91
        40424 => X"53",  -- 83
        40425 => X"51",  -- 81
        40426 => X"59",  -- 89
        40427 => X"55",  -- 85
        40428 => X"4F",  -- 79
        40429 => X"4A",  -- 74
        40430 => X"3C",  -- 60
        40431 => X"39",  -- 57
        40432 => X"2A",  -- 42
        40433 => X"11",  -- 17
        40434 => X"08",  -- 8
        40435 => X"17",  -- 23
        40436 => X"2C",  -- 44
        40437 => X"1F",  -- 31
        40438 => X"8B",  -- 139
        40439 => X"D2",  -- 210
        40440 => X"C2",  -- 194
        40441 => X"B4",  -- 180
        40442 => X"7F",  -- 127
        40443 => X"62",  -- 98
        40444 => X"4B",  -- 75
        40445 => X"40",  -- 64
        40446 => X"58",  -- 88
        40447 => X"5B",  -- 91
        40448 => X"2F",  -- 47
        40449 => X"37",  -- 55
        40450 => X"58",  -- 88
        40451 => X"6F",  -- 111
        40452 => X"69",  -- 105
        40453 => X"62",  -- 98
        40454 => X"72",  -- 114
        40455 => X"84",  -- 132
        40456 => X"8A",  -- 138
        40457 => X"42",  -- 66
        40458 => X"18",  -- 24
        40459 => X"19",  -- 25
        40460 => X"40",  -- 64
        40461 => X"94",  -- 148
        40462 => X"CA",  -- 202
        40463 => X"C6",  -- 198
        40464 => X"D2",  -- 210
        40465 => X"C5",  -- 197
        40466 => X"49",  -- 73
        40467 => X"1B",  -- 27
        40468 => X"76",  -- 118
        40469 => X"C2",  -- 194
        40470 => X"DF",  -- 223
        40471 => X"D5",  -- 213
        40472 => X"D7",  -- 215
        40473 => X"C1",  -- 193
        40474 => X"94",  -- 148
        40475 => X"65",  -- 101
        40476 => X"2C",  -- 44
        40477 => X"18",  -- 24
        40478 => X"2B",  -- 43
        40479 => X"79",  -- 121
        40480 => X"A1",  -- 161
        40481 => X"CB",  -- 203
        40482 => X"CE",  -- 206
        40483 => X"C6",  -- 198
        40484 => X"BE",  -- 190
        40485 => X"AD",  -- 173
        40486 => X"97",  -- 151
        40487 => X"99",  -- 153
        40488 => X"9E",  -- 158
        40489 => X"A9",  -- 169
        40490 => X"C5",  -- 197
        40491 => X"D2",  -- 210
        40492 => X"C7",  -- 199
        40493 => X"BA",  -- 186
        40494 => X"A2",  -- 162
        40495 => X"82",  -- 130
        40496 => X"6E",  -- 110
        40497 => X"72",  -- 114
        40498 => X"73",  -- 115
        40499 => X"6E",  -- 110
        40500 => X"6C",  -- 108
        40501 => X"68",  -- 104
        40502 => X"5D",  -- 93
        40503 => X"50",  -- 80
        40504 => X"63",  -- 99
        40505 => X"55",  -- 85
        40506 => X"46",  -- 70
        40507 => X"3C",  -- 60
        40508 => X"3E",  -- 62
        40509 => X"44",  -- 68
        40510 => X"47",  -- 71
        40511 => X"48",  -- 72
        40512 => X"43",  -- 67
        40513 => X"49",  -- 73
        40514 => X"4F",  -- 79
        40515 => X"55",  -- 85
        40516 => X"5B",  -- 91
        40517 => X"62",  -- 98
        40518 => X"63",  -- 99
        40519 => X"62",  -- 98
        40520 => X"65",  -- 101
        40521 => X"67",  -- 103
        40522 => X"69",  -- 105
        40523 => X"67",  -- 103
        40524 => X"62",  -- 98
        40525 => X"62",  -- 98
        40526 => X"66",  -- 102
        40527 => X"6A",  -- 106
        40528 => X"74",  -- 116
        40529 => X"6E",  -- 110
        40530 => X"67",  -- 103
        40531 => X"65",  -- 101
        40532 => X"68",  -- 104
        40533 => X"6A",  -- 106
        40534 => X"69",  -- 105
        40535 => X"67",  -- 103
        40536 => X"5C",  -- 92
        40537 => X"5D",  -- 93
        40538 => X"61",  -- 97
        40539 => X"60",  -- 96
        40540 => X"57",  -- 87
        40541 => X"4F",  -- 79
        40542 => X"50",  -- 80
        40543 => X"57",  -- 87
        40544 => X"4E",  -- 78
        40545 => X"4D",  -- 77
        40546 => X"46",  -- 70
        40547 => X"40",  -- 64
        40548 => X"40",  -- 64
        40549 => X"44",  -- 68
        40550 => X"46",  -- 70
        40551 => X"45",  -- 69
        40552 => X"48",  -- 72
        40553 => X"5E",  -- 94
        40554 => X"70",  -- 112
        40555 => X"75",  -- 117
        40556 => X"7B",  -- 123
        40557 => X"8A",  -- 138
        40558 => X"9C",  -- 156
        40559 => X"A6",  -- 166
        40560 => X"AF",  -- 175
        40561 => X"BD",  -- 189
        40562 => X"C4",  -- 196
        40563 => X"C1",  -- 193
        40564 => X"C2",  -- 194
        40565 => X"BF",  -- 191
        40566 => X"BA",  -- 186
        40567 => X"BE",  -- 190
        40568 => X"B9",  -- 185
        40569 => X"BD",  -- 189
        40570 => X"B8",  -- 184
        40571 => X"B6",  -- 182
        40572 => X"BA",  -- 186
        40573 => X"B5",  -- 181
        40574 => X"B0",  -- 176
        40575 => X"B6",  -- 182
        40576 => X"A1",  -- 161
        40577 => X"A4",  -- 164
        40578 => X"A4",  -- 164
        40579 => X"B3",  -- 179
        40580 => X"BA",  -- 186
        40581 => X"B2",  -- 178
        40582 => X"B7",  -- 183
        40583 => X"B5",  -- 181
        40584 => X"AA",  -- 170
        40585 => X"A5",  -- 165
        40586 => X"A8",  -- 168
        40587 => X"A8",  -- 168
        40588 => X"AE",  -- 174
        40589 => X"B0",  -- 176
        40590 => X"A5",  -- 165
        40591 => X"AE",  -- 174
        40592 => X"B2",  -- 178
        40593 => X"AB",  -- 171
        40594 => X"A9",  -- 169
        40595 => X"AB",  -- 171
        40596 => X"AD",  -- 173
        40597 => X"B4",  -- 180
        40598 => X"B6",  -- 182
        40599 => X"B0",  -- 176
        40600 => X"B0",  -- 176
        40601 => X"AB",  -- 171
        40602 => X"A3",  -- 163
        40603 => X"A6",  -- 166
        40604 => X"B0",  -- 176
        40605 => X"B3",  -- 179
        40606 => X"B8",  -- 184
        40607 => X"C4",  -- 196
        40608 => X"C7",  -- 199
        40609 => X"C7",  -- 199
        40610 => X"C8",  -- 200
        40611 => X"C9",  -- 201
        40612 => X"C8",  -- 200
        40613 => X"C4",  -- 196
        40614 => X"BE",  -- 190
        40615 => X"B9",  -- 185
        40616 => X"B7",  -- 183
        40617 => X"B6",  -- 182
        40618 => X"B9",  -- 185
        40619 => X"B4",  -- 180
        40620 => X"A4",  -- 164
        40621 => X"94",  -- 148
        40622 => X"8F",  -- 143
        40623 => X"92",  -- 146
        40624 => X"A0",  -- 160
        40625 => X"AD",  -- 173
        40626 => X"A3",  -- 163
        40627 => X"96",  -- 150
        40628 => X"8F",  -- 143
        40629 => X"7A",  -- 122
        40630 => X"72",  -- 114
        40631 => X"89",  -- 137
        40632 => X"A1",  -- 161
        40633 => X"9B",  -- 155
        40634 => X"99",  -- 153
        40635 => X"99",  -- 153
        40636 => X"82",  -- 130
        40637 => X"58",  -- 88
        40638 => X"4D",  -- 77
        40639 => X"67",  -- 103
        40640 => X"4A",  -- 74
        40641 => X"4C",  -- 76
        40642 => X"4D",  -- 77
        40643 => X"4E",  -- 78
        40644 => X"4E",  -- 78
        40645 => X"51",  -- 81
        40646 => X"56",  -- 86
        40647 => X"5B",  -- 91
        40648 => X"58",  -- 88
        40649 => X"58",  -- 88
        40650 => X"55",  -- 85
        40651 => X"4E",  -- 78
        40652 => X"47",  -- 71
        40653 => X"43",  -- 67
        40654 => X"46",  -- 70
        40655 => X"49",  -- 73
        40656 => X"49",  -- 73
        40657 => X"47",  -- 71
        40658 => X"44",  -- 68
        40659 => X"42",  -- 66
        40660 => X"40",  -- 64
        40661 => X"3F",  -- 63
        40662 => X"3D",  -- 61
        40663 => X"3A",  -- 58
        40664 => X"39",  -- 57
        40665 => X"3C",  -- 60
        40666 => X"56",  -- 86
        40667 => X"63",  -- 99
        40668 => X"78",  -- 120
        40669 => X"78",  -- 120
        40670 => X"5E",  -- 94
        40671 => X"6D",  -- 109
        40672 => X"6D",  -- 109
        40673 => X"5E",  -- 94
        40674 => X"48",  -- 72
        40675 => X"33",  -- 51
        40676 => X"13",  -- 19
        40677 => X"08",  -- 8
        40678 => X"21",  -- 33
        40679 => X"34",  -- 52
        40680 => X"82",  -- 130
        40681 => X"9E",  -- 158
        40682 => X"98",  -- 152
        40683 => X"77",  -- 119
        40684 => X"35",  -- 53
        40685 => X"2E",  -- 46
        40686 => X"6A",  -- 106
        40687 => X"81",  -- 129
        40688 => X"71",  -- 113
        40689 => X"62",  -- 98
        40690 => X"1F",  -- 31
        40691 => X"0E",  -- 14
        40692 => X"11",  -- 17
        40693 => X"44",  -- 68
        40694 => X"67",  -- 103
        40695 => X"68",  -- 104
        40696 => X"55",  -- 85
        40697 => X"3E",  -- 62
        40698 => X"3D",  -- 61
        40699 => X"32",  -- 50
        40700 => X"16",  -- 22
        40701 => X"29",  -- 41
        40702 => X"56",  -- 86
        40703 => X"63",  -- 99
        40704 => X"5F",  -- 95
        40705 => X"5D",  -- 93
        40706 => X"4E",  -- 78
        40707 => X"5D",  -- 93
        40708 => X"6C",  -- 108
        40709 => X"92",  -- 146
        40710 => X"A7",  -- 167
        40711 => X"64",  -- 100
        40712 => X"09",  -- 9
        40713 => X"0F",  -- 15
        40714 => X"06",  -- 6
        40715 => X"12",  -- 18
        40716 => X"11",  -- 17
        40717 => X"1E",  -- 30
        40718 => X"14",  -- 20
        40719 => X"1E",  -- 30
        40720 => X"22",  -- 34
        40721 => X"27",  -- 39
        40722 => X"2D",  -- 45
        40723 => X"2E",  -- 46
        40724 => X"2E",  -- 46
        40725 => X"30",  -- 48
        40726 => X"37",  -- 55
        40727 => X"3C",  -- 60
        40728 => X"43",  -- 67
        40729 => X"50",  -- 80
        40730 => X"58",  -- 88
        40731 => X"54",  -- 84
        40732 => X"64",  -- 100
        40733 => X"49",  -- 73
        40734 => X"4D",  -- 77
        40735 => X"6B",  -- 107
        40736 => X"68",  -- 104
        40737 => X"67",  -- 103
        40738 => X"5B",  -- 91
        40739 => X"63",  -- 99
        40740 => X"69",  -- 105
        40741 => X"5E",  -- 94
        40742 => X"64",  -- 100
        40743 => X"6C",  -- 108
        40744 => X"59",  -- 89
        40745 => X"57",  -- 87
        40746 => X"69",  -- 105
        40747 => X"5D",  -- 93
        40748 => X"51",  -- 81
        40749 => X"4B",  -- 75
        40750 => X"34",  -- 52
        40751 => X"36",  -- 54
        40752 => X"30",  -- 48
        40753 => X"15",  -- 21
        40754 => X"18",  -- 24
        40755 => X"16",  -- 22
        40756 => X"1A",  -- 26
        40757 => X"29",  -- 41
        40758 => X"9D",  -- 157
        40759 => X"CB",  -- 203
        40760 => X"B6",  -- 182
        40761 => X"93",  -- 147
        40762 => X"83",  -- 131
        40763 => X"62",  -- 98
        40764 => X"5A",  -- 90
        40765 => X"6B",  -- 107
        40766 => X"61",  -- 97
        40767 => X"63",  -- 99
        40768 => X"48",  -- 72
        40769 => X"4E",  -- 78
        40770 => X"67",  -- 103
        40771 => X"80",  -- 128
        40772 => X"83",  -- 131
        40773 => X"82",  -- 130
        40774 => X"89",  -- 137
        40775 => X"8F",  -- 143
        40776 => X"66",  -- 102
        40777 => X"39",  -- 57
        40778 => X"18",  -- 24
        40779 => X"14",  -- 20
        40780 => X"43",  -- 67
        40781 => X"A6",  -- 166
        40782 => X"CB",  -- 203
        40783 => X"B0",  -- 176
        40784 => X"CD",  -- 205
        40785 => X"C4",  -- 196
        40786 => X"4C",  -- 76
        40787 => X"27",  -- 39
        40788 => X"85",  -- 133
        40789 => X"C8",  -- 200
        40790 => X"E1",  -- 225
        40791 => X"D6",  -- 214
        40792 => X"D3",  -- 211
        40793 => X"C6",  -- 198
        40794 => X"9C",  -- 156
        40795 => X"73",  -- 115
        40796 => X"3C",  -- 60
        40797 => X"1E",  -- 30
        40798 => X"21",  -- 33
        40799 => X"69",  -- 105
        40800 => X"9A",  -- 154
        40801 => X"C7",  -- 199
        40802 => X"D1",  -- 209
        40803 => X"CA",  -- 202
        40804 => X"C0",  -- 192
        40805 => X"BC",  -- 188
        40806 => X"93",  -- 147
        40807 => X"91",  -- 145
        40808 => X"AC",  -- 172
        40809 => X"A4",  -- 164
        40810 => X"BE",  -- 190
        40811 => X"D7",  -- 215
        40812 => X"C3",  -- 195
        40813 => X"AE",  -- 174
        40814 => X"A4",  -- 164
        40815 => X"96",  -- 150
        40816 => X"79",  -- 121
        40817 => X"7F",  -- 127
        40818 => X"7D",  -- 125
        40819 => X"76",  -- 118
        40820 => X"73",  -- 115
        40821 => X"6E",  -- 110
        40822 => X"5A",  -- 90
        40823 => X"43",  -- 67
        40824 => X"4A",  -- 74
        40825 => X"50",  -- 80
        40826 => X"57",  -- 87
        40827 => X"55",  -- 85
        40828 => X"4A",  -- 74
        40829 => X"40",  -- 64
        40830 => X"3E",  -- 62
        40831 => X"44",  -- 68
        40832 => X"4B",  -- 75
        40833 => X"4D",  -- 77
        40834 => X"4F",  -- 79
        40835 => X"50",  -- 80
        40836 => X"5A",  -- 90
        40837 => X"66",  -- 102
        40838 => X"6B",  -- 107
        40839 => X"68",  -- 104
        40840 => X"61",  -- 97
        40841 => X"66",  -- 102
        40842 => X"6B",  -- 107
        40843 => X"69",  -- 105
        40844 => X"62",  -- 98
        40845 => X"5E",  -- 94
        40846 => X"60",  -- 96
        40847 => X"63",  -- 99
        40848 => X"6D",  -- 109
        40849 => X"69",  -- 105
        40850 => X"65",  -- 101
        40851 => X"63",  -- 99
        40852 => X"63",  -- 99
        40853 => X"63",  -- 99
        40854 => X"61",  -- 97
        40855 => X"5F",  -- 95
        40856 => X"5C",  -- 92
        40857 => X"57",  -- 87
        40858 => X"55",  -- 85
        40859 => X"59",  -- 89
        40860 => X"5A",  -- 90
        40861 => X"54",  -- 84
        40862 => X"4D",  -- 77
        40863 => X"4C",  -- 76
        40864 => X"4F",  -- 79
        40865 => X"4C",  -- 76
        40866 => X"45",  -- 69
        40867 => X"3E",  -- 62
        40868 => X"3D",  -- 61
        40869 => X"42",  -- 66
        40870 => X"45",  -- 69
        40871 => X"45",  -- 69
        40872 => X"54",  -- 84
        40873 => X"69",  -- 105
        40874 => X"78",  -- 120
        40875 => X"7B",  -- 123
        40876 => X"7E",  -- 126
        40877 => X"8E",  -- 142
        40878 => X"A1",  -- 161
        40879 => X"AC",  -- 172
        40880 => X"A9",  -- 169
        40881 => X"B8",  -- 184
        40882 => X"C2",  -- 194
        40883 => X"C5",  -- 197
        40884 => X"C6",  -- 198
        40885 => X"BD",  -- 189
        40886 => X"B9",  -- 185
        40887 => X"C1",  -- 193
        40888 => X"B8",  -- 184
        40889 => X"B6",  -- 182
        40890 => X"B1",  -- 177
        40891 => X"AF",  -- 175
        40892 => X"B1",  -- 177
        40893 => X"AB",  -- 171
        40894 => X"AB",  -- 171
        40895 => X"B7",  -- 183
        40896 => X"A0",  -- 160
        40897 => X"A0",  -- 160
        40898 => X"A1",  -- 161
        40899 => X"B3",  -- 179
        40900 => X"B9",  -- 185
        40901 => X"AE",  -- 174
        40902 => X"B3",  -- 179
        40903 => X"B3",  -- 179
        40904 => X"A5",  -- 165
        40905 => X"A2",  -- 162
        40906 => X"A6",  -- 166
        40907 => X"A3",  -- 163
        40908 => X"AF",  -- 175
        40909 => X"B2",  -- 178
        40910 => X"A6",  -- 166
        40911 => X"AB",  -- 171
        40912 => X"BA",  -- 186
        40913 => X"A8",  -- 168
        40914 => X"A9",  -- 169
        40915 => X"B0",  -- 176
        40916 => X"B0",  -- 176
        40917 => X"B5",  -- 181
        40918 => X"B8",  -- 184
        40919 => X"AD",  -- 173
        40920 => X"AA",  -- 170
        40921 => X"B4",  -- 180
        40922 => X"AB",  -- 171
        40923 => X"A4",  -- 164
        40924 => X"B0",  -- 176
        40925 => X"B6",  -- 182
        40926 => X"BA",  -- 186
        40927 => X"C6",  -- 198
        40928 => X"CA",  -- 202
        40929 => X"C8",  -- 200
        40930 => X"C8",  -- 200
        40931 => X"C8",  -- 200
        40932 => X"C8",  -- 200
        40933 => X"C4",  -- 196
        40934 => X"BC",  -- 188
        40935 => X"B5",  -- 181
        40936 => X"B0",  -- 176
        40937 => X"B6",  -- 182
        40938 => X"BB",  -- 187
        40939 => X"BB",  -- 187
        40940 => X"B2",  -- 178
        40941 => X"A5",  -- 165
        40942 => X"98",  -- 152
        40943 => X"90",  -- 144
        40944 => X"94",  -- 148
        40945 => X"AB",  -- 171
        40946 => X"9F",  -- 159
        40947 => X"88",  -- 136
        40948 => X"84",  -- 132
        40949 => X"79",  -- 121
        40950 => X"6D",  -- 109
        40951 => X"75",  -- 117
        40952 => X"96",  -- 150
        40953 => X"AD",  -- 173
        40954 => X"99",  -- 153
        40955 => X"85",  -- 133
        40956 => X"8B",  -- 139
        40957 => X"6A",  -- 106
        40958 => X"48",  -- 72
        40959 => X"59",  -- 89
        40960 => X"4D",  -- 77
        40961 => X"4E",  -- 78
        40962 => X"51",  -- 81
        40963 => X"55",  -- 85
        40964 => X"58",  -- 88
        40965 => X"5C",  -- 92
        40966 => X"60",  -- 96
        40967 => X"63",  -- 99
        40968 => X"60",  -- 96
        40969 => X"5E",  -- 94
        40970 => X"59",  -- 89
        40971 => X"53",  -- 83
        40972 => X"4E",  -- 78
        40973 => X"4A",  -- 74
        40974 => X"46",  -- 70
        40975 => X"45",  -- 69
        40976 => X"44",  -- 68
        40977 => X"46",  -- 70
        40978 => X"48",  -- 72
        40979 => X"47",  -- 71
        40980 => X"45",  -- 69
        40981 => X"41",  -- 65
        40982 => X"3C",  -- 60
        40983 => X"3C",  -- 60
        40984 => X"3C",  -- 60
        40985 => X"3F",  -- 63
        40986 => X"5A",  -- 90
        40987 => X"6E",  -- 110
        40988 => X"65",  -- 101
        40989 => X"63",  -- 99
        40990 => X"71",  -- 113
        40991 => X"75",  -- 117
        40992 => X"64",  -- 100
        40993 => X"5C",  -- 92
        40994 => X"56",  -- 86
        40995 => X"34",  -- 52
        40996 => X"14",  -- 20
        40997 => X"0B",  -- 11
        40998 => X"17",  -- 23
        40999 => X"39",  -- 57
        41000 => X"8E",  -- 142
        41001 => X"9B",  -- 155
        41002 => X"96",  -- 150
        41003 => X"89",  -- 137
        41004 => X"4A",  -- 74
        41005 => X"1B",  -- 27
        41006 => X"51",  -- 81
        41007 => X"8D",  -- 141
        41008 => X"72",  -- 114
        41009 => X"68",  -- 104
        41010 => X"44",  -- 68
        41011 => X"07",  -- 7
        41012 => X"0A",  -- 10
        41013 => X"31",  -- 49
        41014 => X"3E",  -- 62
        41015 => X"5B",  -- 91
        41016 => X"4E",  -- 78
        41017 => X"65",  -- 101
        41018 => X"5F",  -- 95
        41019 => X"3F",  -- 63
        41020 => X"3A",  -- 58
        41021 => X"4C",  -- 76
        41022 => X"51",  -- 81
        41023 => X"4C",  -- 76
        41024 => X"42",  -- 66
        41025 => X"51",  -- 81
        41026 => X"4D",  -- 77
        41027 => X"5F",  -- 95
        41028 => X"6D",  -- 109
        41029 => X"84",  -- 132
        41030 => X"8D",  -- 141
        41031 => X"45",  -- 69
        41032 => X"17",  -- 23
        41033 => X"1E",  -- 30
        41034 => X"1A",  -- 26
        41035 => X"14",  -- 20
        41036 => X"1F",  -- 31
        41037 => X"26",  -- 38
        41038 => X"21",  -- 33
        41039 => X"1D",  -- 29
        41040 => X"27",  -- 39
        41041 => X"26",  -- 38
        41042 => X"2A",  -- 42
        41043 => X"2F",  -- 47
        41044 => X"31",  -- 49
        41045 => X"33",  -- 51
        41046 => X"36",  -- 54
        41047 => X"3C",  -- 60
        41048 => X"4D",  -- 77
        41049 => X"4B",  -- 75
        41050 => X"54",  -- 84
        41051 => X"61",  -- 97
        41052 => X"60",  -- 96
        41053 => X"56",  -- 86
        41054 => X"57",  -- 87
        41055 => X"60",  -- 96
        41056 => X"65",  -- 101
        41057 => X"70",  -- 112
        41058 => X"6C",  -- 108
        41059 => X"75",  -- 117
        41060 => X"6C",  -- 108
        41061 => X"6B",  -- 107
        41062 => X"60",  -- 96
        41063 => X"6A",  -- 106
        41064 => X"5E",  -- 94
        41065 => X"55",  -- 85
        41066 => X"59",  -- 89
        41067 => X"65",  -- 101
        41068 => X"5F",  -- 95
        41069 => X"48",  -- 72
        41070 => X"3D",  -- 61
        41071 => X"40",  -- 64
        41072 => X"3F",  -- 63
        41073 => X"33",  -- 51
        41074 => X"0E",  -- 14
        41075 => X"1A",  -- 26
        41076 => X"1D",  -- 29
        41077 => X"30",  -- 48
        41078 => X"94",  -- 148
        41079 => X"C5",  -- 197
        41080 => X"9B",  -- 155
        41081 => X"85",  -- 133
        41082 => X"77",  -- 119
        41083 => X"72",  -- 114
        41084 => X"6B",  -- 107
        41085 => X"6B",  -- 107
        41086 => X"70",  -- 112
        41087 => X"6C",  -- 108
        41088 => X"69",  -- 105
        41089 => X"71",  -- 113
        41090 => X"79",  -- 121
        41091 => X"89",  -- 137
        41092 => X"8F",  -- 143
        41093 => X"8B",  -- 139
        41094 => X"88",  -- 136
        41095 => X"82",  -- 130
        41096 => X"77",  -- 119
        41097 => X"37",  -- 55
        41098 => X"16",  -- 22
        41099 => X"1B",  -- 27
        41100 => X"5C",  -- 92
        41101 => X"B2",  -- 178
        41102 => X"BA",  -- 186
        41103 => X"A0",  -- 160
        41104 => X"CF",  -- 207
        41105 => X"C5",  -- 197
        41106 => X"42",  -- 66
        41107 => X"3F",  -- 63
        41108 => X"98",  -- 152
        41109 => X"CF",  -- 207
        41110 => X"D7",  -- 215
        41111 => X"D9",  -- 217
        41112 => X"D2",  -- 210
        41113 => X"CC",  -- 204
        41114 => X"99",  -- 153
        41115 => X"5C",  -- 92
        41116 => X"48",  -- 72
        41117 => X"1E",  -- 30
        41118 => X"17",  -- 23
        41119 => X"57",  -- 87
        41120 => X"99",  -- 153
        41121 => X"BB",  -- 187
        41122 => X"D1",  -- 209
        41123 => X"CD",  -- 205
        41124 => X"B8",  -- 184
        41125 => X"B8",  -- 184
        41126 => X"B0",  -- 176
        41127 => X"7C",  -- 124
        41128 => X"9D",  -- 157
        41129 => X"B9",  -- 185
        41130 => X"B7",  -- 183
        41131 => X"CE",  -- 206
        41132 => X"D6",  -- 214
        41133 => X"9C",  -- 156
        41134 => X"81",  -- 129
        41135 => X"9F",  -- 159
        41136 => X"87",  -- 135
        41137 => X"74",  -- 116
        41138 => X"81",  -- 129
        41139 => X"77",  -- 119
        41140 => X"70",  -- 112
        41141 => X"7A",  -- 122
        41142 => X"64",  -- 100
        41143 => X"52",  -- 82
        41144 => X"49",  -- 73
        41145 => X"4A",  -- 74
        41146 => X"4C",  -- 76
        41147 => X"52",  -- 82
        41148 => X"56",  -- 86
        41149 => X"54",  -- 84
        41150 => X"4E",  -- 78
        41151 => X"48",  -- 72
        41152 => X"51",  -- 81
        41153 => X"56",  -- 86
        41154 => X"59",  -- 89
        41155 => X"58",  -- 88
        41156 => X"5B",  -- 91
        41157 => X"62",  -- 98
        41158 => X"66",  -- 102
        41159 => X"65",  -- 101
        41160 => X"6A",  -- 106
        41161 => X"67",  -- 103
        41162 => X"68",  -- 104
        41163 => X"66",  -- 102
        41164 => X"5D",  -- 93
        41165 => X"55",  -- 85
        41166 => X"5C",  -- 92
        41167 => X"6A",  -- 106
        41168 => X"65",  -- 101
        41169 => X"65",  -- 101
        41170 => X"61",  -- 97
        41171 => X"5D",  -- 93
        41172 => X"5E",  -- 94
        41173 => X"61",  -- 97
        41174 => X"5D",  -- 93
        41175 => X"56",  -- 86
        41176 => X"53",  -- 83
        41177 => X"54",  -- 84
        41178 => X"56",  -- 86
        41179 => X"55",  -- 85
        41180 => X"52",  -- 82
        41181 => X"4E",  -- 78
        41182 => X"4C",  -- 76
        41183 => X"4B",  -- 75
        41184 => X"49",  -- 73
        41185 => X"4C",  -- 76
        41186 => X"46",  -- 70
        41187 => X"3E",  -- 62
        41188 => X"42",  -- 66
        41189 => X"41",  -- 65
        41190 => X"42",  -- 66
        41191 => X"4A",  -- 74
        41192 => X"61",  -- 97
        41193 => X"6D",  -- 109
        41194 => X"77",  -- 119
        41195 => X"7D",  -- 125
        41196 => X"86",  -- 134
        41197 => X"97",  -- 151
        41198 => X"A7",  -- 167
        41199 => X"B2",  -- 178
        41200 => X"B4",  -- 180
        41201 => X"BB",  -- 187
        41202 => X"CD",  -- 205
        41203 => X"CB",  -- 203
        41204 => X"C5",  -- 197
        41205 => X"C4",  -- 196
        41206 => X"BC",  -- 188
        41207 => X"BF",  -- 191
        41208 => X"BC",  -- 188
        41209 => X"B9",  -- 185
        41210 => X"B3",  -- 179
        41211 => X"B1",  -- 177
        41212 => X"B0",  -- 176
        41213 => X"A7",  -- 167
        41214 => X"A6",  -- 166
        41215 => X"B2",  -- 178
        41216 => X"97",  -- 151
        41217 => X"A1",  -- 161
        41218 => X"A4",  -- 164
        41219 => X"AA",  -- 170
        41220 => X"B7",  -- 183
        41221 => X"AE",  -- 174
        41222 => X"A4",  -- 164
        41223 => X"AF",  -- 175
        41224 => X"9F",  -- 159
        41225 => X"9E",  -- 158
        41226 => X"9E",  -- 158
        41227 => X"A4",  -- 164
        41228 => X"A9",  -- 169
        41229 => X"AD",  -- 173
        41230 => X"AB",  -- 171
        41231 => X"A9",  -- 169
        41232 => X"B2",  -- 178
        41233 => X"B3",  -- 179
        41234 => X"AE",  -- 174
        41235 => X"A8",  -- 168
        41236 => X"AA",  -- 170
        41237 => X"B2",  -- 178
        41238 => X"B4",  -- 180
        41239 => X"B0",  -- 176
        41240 => X"AF",  -- 175
        41241 => X"AA",  -- 170
        41242 => X"A9",  -- 169
        41243 => X"AB",  -- 171
        41244 => X"AC",  -- 172
        41245 => X"B1",  -- 177
        41246 => X"BB",  -- 187
        41247 => X"C5",  -- 197
        41248 => X"C8",  -- 200
        41249 => X"CA",  -- 202
        41250 => X"CB",  -- 203
        41251 => X"CB",  -- 203
        41252 => X"CC",  -- 204
        41253 => X"C7",  -- 199
        41254 => X"B9",  -- 185
        41255 => X"AB",  -- 171
        41256 => X"A3",  -- 163
        41257 => X"A6",  -- 166
        41258 => X"B5",  -- 181
        41259 => X"BF",  -- 191
        41260 => X"B9",  -- 185
        41261 => X"B1",  -- 177
        41262 => X"A8",  -- 168
        41263 => X"99",  -- 153
        41264 => X"A1",  -- 161
        41265 => X"9F",  -- 159
        41266 => X"9A",  -- 154
        41267 => X"A4",  -- 164
        41268 => X"82",  -- 130
        41269 => X"5B",  -- 91
        41270 => X"6A",  -- 106
        41271 => X"65",  -- 101
        41272 => X"88",  -- 136
        41273 => X"9F",  -- 159
        41274 => X"AA",  -- 170
        41275 => X"97",  -- 151
        41276 => X"7B",  -- 123
        41277 => X"6A",  -- 106
        41278 => X"5A",  -- 90
        41279 => X"4E",  -- 78
        41280 => X"57",  -- 87
        41281 => X"55",  -- 85
        41282 => X"56",  -- 86
        41283 => X"5A",  -- 90
        41284 => X"63",  -- 99
        41285 => X"6C",  -- 108
        41286 => X"70",  -- 112
        41287 => X"71",  -- 113
        41288 => X"6E",  -- 110
        41289 => X"6A",  -- 106
        41290 => X"65",  -- 101
        41291 => X"5F",  -- 95
        41292 => X"58",  -- 88
        41293 => X"52",  -- 82
        41294 => X"4D",  -- 77
        41295 => X"4B",  -- 75
        41296 => X"45",  -- 69
        41297 => X"46",  -- 70
        41298 => X"49",  -- 73
        41299 => X"48",  -- 72
        41300 => X"46",  -- 70
        41301 => X"44",  -- 68
        41302 => X"43",  -- 67
        41303 => X"43",  -- 67
        41304 => X"46",  -- 70
        41305 => X"47",  -- 71
        41306 => X"5A",  -- 90
        41307 => X"68",  -- 104
        41308 => X"62",  -- 98
        41309 => X"64",  -- 100
        41310 => X"68",  -- 104
        41311 => X"64",  -- 100
        41312 => X"61",  -- 97
        41313 => X"62",  -- 98
        41314 => X"59",  -- 89
        41315 => X"33",  -- 51
        41316 => X"18",  -- 24
        41317 => X"12",  -- 18
        41318 => X"1F",  -- 31
        41319 => X"47",  -- 71
        41320 => X"90",  -- 144
        41321 => X"A0",  -- 160
        41322 => X"97",  -- 151
        41323 => X"8D",  -- 141
        41324 => X"68",  -- 104
        41325 => X"26",  -- 38
        41326 => X"35",  -- 53
        41327 => X"7E",  -- 126
        41328 => X"8E",  -- 142
        41329 => X"76",  -- 118
        41330 => X"56",  -- 86
        41331 => X"1F",  -- 31
        41332 => X"04",  -- 4
        41333 => X"18",  -- 24
        41334 => X"22",  -- 34
        41335 => X"1A",  -- 26
        41336 => X"3B",  -- 59
        41337 => X"4D",  -- 77
        41338 => X"5B",  -- 91
        41339 => X"61",  -- 97
        41340 => X"62",  -- 98
        41341 => X"57",  -- 87
        41342 => X"50",  -- 80
        41343 => X"52",  -- 82
        41344 => X"49",  -- 73
        41345 => X"5E",  -- 94
        41346 => X"5E",  -- 94
        41347 => X"66",  -- 102
        41348 => X"64",  -- 100
        41349 => X"6F",  -- 111
        41350 => X"7E",  -- 126
        41351 => X"49",  -- 73
        41352 => X"30",  -- 48
        41353 => X"2A",  -- 42
        41354 => X"1C",  -- 28
        41355 => X"19",  -- 25
        41356 => X"26",  -- 38
        41357 => X"2A",  -- 42
        41358 => X"23",  -- 35
        41359 => X"1E",  -- 30
        41360 => X"29",  -- 41
        41361 => X"29",  -- 41
        41362 => X"2B",  -- 43
        41363 => X"30",  -- 48
        41364 => X"34",  -- 52
        41365 => X"38",  -- 56
        41366 => X"3D",  -- 61
        41367 => X"44",  -- 68
        41368 => X"4D",  -- 77
        41369 => X"4E",  -- 78
        41370 => X"50",  -- 80
        41371 => X"52",  -- 82
        41372 => X"53",  -- 83
        41373 => X"57",  -- 87
        41374 => X"60",  -- 96
        41375 => X"67",  -- 103
        41376 => X"6B",  -- 107
        41377 => X"77",  -- 119
        41378 => X"6C",  -- 108
        41379 => X"6B",  -- 107
        41380 => X"63",  -- 99
        41381 => X"69",  -- 105
        41382 => X"5C",  -- 92
        41383 => X"5E",  -- 94
        41384 => X"69",  -- 105
        41385 => X"60",  -- 96
        41386 => X"5E",  -- 94
        41387 => X"62",  -- 98
        41388 => X"5C",  -- 92
        41389 => X"4C",  -- 76
        41390 => X"44",  -- 68
        41391 => X"47",  -- 71
        41392 => X"46",  -- 70
        41393 => X"32",  -- 50
        41394 => X"1A",  -- 26
        41395 => X"30",  -- 48
        41396 => X"3F",  -- 63
        41397 => X"4F",  -- 79
        41398 => X"89",  -- 137
        41399 => X"A4",  -- 164
        41400 => X"90",  -- 144
        41401 => X"7D",  -- 125
        41402 => X"72",  -- 114
        41403 => X"6E",  -- 110
        41404 => X"67",  -- 103
        41405 => X"65",  -- 101
        41406 => X"65",  -- 101
        41407 => X"60",  -- 96
        41408 => X"6F",  -- 111
        41409 => X"78",  -- 120
        41410 => X"76",  -- 118
        41411 => X"76",  -- 118
        41412 => X"7A",  -- 122
        41413 => X"83",  -- 131
        41414 => X"8E",  -- 142
        41415 => X"91",  -- 145
        41416 => X"8C",  -- 140
        41417 => X"30",  -- 48
        41418 => X"02",  -- 2
        41419 => X"26",  -- 38
        41420 => X"84",  -- 132
        41421 => X"CD",  -- 205
        41422 => X"C9",  -- 201
        41423 => X"B5",  -- 181
        41424 => X"D0",  -- 208
        41425 => X"B8",  -- 184
        41426 => X"50",  -- 80
        41427 => X"60",  -- 96
        41428 => X"AB",  -- 171
        41429 => X"CE",  -- 206
        41430 => X"D1",  -- 209
        41431 => X"D5",  -- 213
        41432 => X"D3",  -- 211
        41433 => X"CB",  -- 203
        41434 => X"99",  -- 153
        41435 => X"51",  -- 81
        41436 => X"3C",  -- 60
        41437 => X"2A",  -- 42
        41438 => X"1A",  -- 26
        41439 => X"47",  -- 71
        41440 => X"8B",  -- 139
        41441 => X"BF",  -- 191
        41442 => X"D4",  -- 212
        41443 => X"C7",  -- 199
        41444 => X"B4",  -- 180
        41445 => X"AB",  -- 171
        41446 => X"AB",  -- 171
        41447 => X"9D",  -- 157
        41448 => X"A1",  -- 161
        41449 => X"AE",  -- 174
        41450 => X"B9",  -- 185
        41451 => X"C9",  -- 201
        41452 => X"D7",  -- 215
        41453 => X"B3",  -- 179
        41454 => X"7E",  -- 126
        41455 => X"81",  -- 129
        41456 => X"89",  -- 137
        41457 => X"7D",  -- 125
        41458 => X"73",  -- 115
        41459 => X"75",  -- 117
        41460 => X"73",  -- 115
        41461 => X"6E",  -- 110
        41462 => X"6B",  -- 107
        41463 => X"60",  -- 96
        41464 => X"5A",  -- 90
        41465 => X"54",  -- 84
        41466 => X"4E",  -- 78
        41467 => X"4D",  -- 77
        41468 => X"50",  -- 80
        41469 => X"54",  -- 84
        41470 => X"53",  -- 83
        41471 => X"51",  -- 81
        41472 => X"55",  -- 85
        41473 => X"59",  -- 89
        41474 => X"5B",  -- 91
        41475 => X"59",  -- 89
        41476 => X"5A",  -- 90
        41477 => X"60",  -- 96
        41478 => X"64",  -- 100
        41479 => X"65",  -- 101
        41480 => X"65",  -- 101
        41481 => X"63",  -- 99
        41482 => X"65",  -- 101
        41483 => X"66",  -- 102
        41484 => X"5F",  -- 95
        41485 => X"57",  -- 87
        41486 => X"59",  -- 89
        41487 => X"63",  -- 99
        41488 => X"63",  -- 99
        41489 => X"62",  -- 98
        41490 => X"5E",  -- 94
        41491 => X"5A",  -- 90
        41492 => X"5B",  -- 91
        41493 => X"5D",  -- 93
        41494 => X"5A",  -- 90
        41495 => X"54",  -- 84
        41496 => X"4D",  -- 77
        41497 => X"50",  -- 80
        41498 => X"53",  -- 83
        41499 => X"54",  -- 84
        41500 => X"51",  -- 81
        41501 => X"4D",  -- 77
        41502 => X"49",  -- 73
        41503 => X"48",  -- 72
        41504 => X"48",  -- 72
        41505 => X"4C",  -- 76
        41506 => X"45",  -- 69
        41507 => X"3F",  -- 63
        41508 => X"42",  -- 66
        41509 => X"42",  -- 66
        41510 => X"45",  -- 69
        41511 => X"4C",  -- 76
        41512 => X"66",  -- 102
        41513 => X"6F",  -- 111
        41514 => X"7B",  -- 123
        41515 => X"81",  -- 129
        41516 => X"8C",  -- 140
        41517 => X"9E",  -- 158
        41518 => X"AC",  -- 172
        41519 => X"B5",  -- 181
        41520 => X"BC",  -- 188
        41521 => X"BF",  -- 191
        41522 => X"CB",  -- 203
        41523 => X"C8",  -- 200
        41524 => X"C7",  -- 199
        41525 => X"C9",  -- 201
        41526 => X"BD",  -- 189
        41527 => X"BB",  -- 187
        41528 => X"C5",  -- 197
        41529 => X"C0",  -- 192
        41530 => X"B9",  -- 185
        41531 => X"B3",  -- 179
        41532 => X"AA",  -- 170
        41533 => X"A4",  -- 164
        41534 => X"A5",  -- 165
        41535 => X"A8",  -- 168
        41536 => X"97",  -- 151
        41537 => X"9A",  -- 154
        41538 => X"9F",  -- 159
        41539 => X"A7",  -- 167
        41540 => X"AB",  -- 171
        41541 => X"A3",  -- 163
        41542 => X"A1",  -- 161
        41543 => X"AA",  -- 170
        41544 => X"A1",  -- 161
        41545 => X"9F",  -- 159
        41546 => X"9D",  -- 157
        41547 => X"9D",  -- 157
        41548 => X"9E",  -- 158
        41549 => X"9F",  -- 159
        41550 => X"A1",  -- 161
        41551 => X"A1",  -- 161
        41552 => X"AE",  -- 174
        41553 => X"B3",  -- 179
        41554 => X"B2",  -- 178
        41555 => X"AB",  -- 171
        41556 => X"A9",  -- 169
        41557 => X"AF",  -- 175
        41558 => X"B2",  -- 178
        41559 => X"B0",  -- 176
        41560 => X"AC",  -- 172
        41561 => X"AA",  -- 170
        41562 => X"AA",  -- 170
        41563 => X"AD",  -- 173
        41564 => X"AF",  -- 175
        41565 => X"B2",  -- 178
        41566 => X"BC",  -- 188
        41567 => X"C6",  -- 198
        41568 => X"C8",  -- 200
        41569 => X"CB",  -- 203
        41570 => X"CA",  -- 202
        41571 => X"C9",  -- 201
        41572 => X"C8",  -- 200
        41573 => X"C4",  -- 196
        41574 => X"BA",  -- 186
        41575 => X"AF",  -- 175
        41576 => X"A0",  -- 160
        41577 => X"9D",  -- 157
        41578 => X"A6",  -- 166
        41579 => X"B1",  -- 177
        41580 => X"B3",  -- 179
        41581 => X"B3",  -- 179
        41582 => X"AC",  -- 172
        41583 => X"9F",  -- 159
        41584 => X"98",  -- 152
        41585 => X"A0",  -- 160
        41586 => X"A0",  -- 160
        41587 => X"88",  -- 136
        41588 => X"87",  -- 135
        41589 => X"75",  -- 117
        41590 => X"4C",  -- 76
        41591 => X"5F",  -- 95
        41592 => X"77",  -- 119
        41593 => X"8F",  -- 143
        41594 => X"A5",  -- 165
        41595 => X"9E",  -- 158
        41596 => X"84",  -- 132
        41597 => X"68",  -- 104
        41598 => X"58",  -- 88
        41599 => X"53",  -- 83
        41600 => X"61",  -- 97
        41601 => X"5D",  -- 93
        41602 => X"5B",  -- 91
        41603 => X"5F",  -- 95
        41604 => X"6C",  -- 108
        41605 => X"7B",  -- 123
        41606 => X"82",  -- 130
        41607 => X"85",  -- 133
        41608 => X"83",  -- 131
        41609 => X"7E",  -- 126
        41610 => X"76",  -- 118
        41611 => X"6F",  -- 111
        41612 => X"69",  -- 105
        41613 => X"61",  -- 97
        41614 => X"58",  -- 88
        41615 => X"51",  -- 81
        41616 => X"4B",  -- 75
        41617 => X"4A",  -- 74
        41618 => X"4A",  -- 74
        41619 => X"49",  -- 73
        41620 => X"49",  -- 73
        41621 => X"4B",  -- 75
        41622 => X"4B",  -- 75
        41623 => X"4C",  -- 76
        41624 => X"4F",  -- 79
        41625 => X"4F",  -- 79
        41626 => X"5A",  -- 90
        41627 => X"62",  -- 98
        41628 => X"64",  -- 100
        41629 => X"66",  -- 102
        41630 => X"62",  -- 98
        41631 => X"52",  -- 82
        41632 => X"58",  -- 88
        41633 => X"66",  -- 102
        41634 => X"5A",  -- 90
        41635 => X"2C",  -- 44
        41636 => X"17",  -- 23
        41637 => X"12",  -- 18
        41638 => X"1D",  -- 29
        41639 => X"4B",  -- 75
        41640 => X"89",  -- 137
        41641 => X"97",  -- 151
        41642 => X"8F",  -- 143
        41643 => X"88",  -- 136
        41644 => X"7D",  -- 125
        41645 => X"33",  -- 51
        41646 => X"19",  -- 25
        41647 => X"6C",  -- 108
        41648 => X"8A",  -- 138
        41649 => X"85",  -- 133
        41650 => X"71",  -- 113
        41651 => X"3D",  -- 61
        41652 => X"07",  -- 7
        41653 => X"1F",  -- 31
        41654 => X"3B",  -- 59
        41655 => X"11",  -- 17
        41656 => X"1C",  -- 28
        41657 => X"44",  -- 68
        41658 => X"61",  -- 97
        41659 => X"67",  -- 103
        41660 => X"6E",  -- 110
        41661 => X"6D",  -- 109
        41662 => X"62",  -- 98
        41663 => X"5A",  -- 90
        41664 => X"54",  -- 84
        41665 => X"64",  -- 100
        41666 => X"63",  -- 99
        41667 => X"6A",  -- 106
        41668 => X"61",  -- 97
        41669 => X"62",  -- 98
        41670 => X"70",  -- 112
        41671 => X"4E",  -- 78
        41672 => X"37",  -- 55
        41673 => X"2A",  -- 42
        41674 => X"18",  -- 24
        41675 => X"20",  -- 32
        41676 => X"35",  -- 53
        41677 => X"39",  -- 57
        41678 => X"2D",  -- 45
        41679 => X"28",  -- 40
        41680 => X"2C",  -- 44
        41681 => X"2B",  -- 43
        41682 => X"2F",  -- 47
        41683 => X"34",  -- 52
        41684 => X"39",  -- 57
        41685 => X"3C",  -- 60
        41686 => X"44",  -- 68
        41687 => X"4A",  -- 74
        41688 => X"4F",  -- 79
        41689 => X"56",  -- 86
        41690 => X"58",  -- 88
        41691 => X"52",  -- 82
        41692 => X"4E",  -- 78
        41693 => X"50",  -- 80
        41694 => X"4E",  -- 78
        41695 => X"4B",  -- 75
        41696 => X"57",  -- 87
        41697 => X"68",  -- 104
        41698 => X"62",  -- 98
        41699 => X"65",  -- 101
        41700 => X"68",  -- 104
        41701 => X"78",  -- 120
        41702 => X"6C",  -- 108
        41703 => X"67",  -- 103
        41704 => X"68",  -- 104
        41705 => X"62",  -- 98
        41706 => X"5D",  -- 93
        41707 => X"58",  -- 88
        41708 => X"53",  -- 83
        41709 => X"4E",  -- 78
        41710 => X"4D",  -- 77
        41711 => X"4D",  -- 77
        41712 => X"4C",  -- 76
        41713 => X"2B",  -- 43
        41714 => X"1D",  -- 29
        41715 => X"2A",  -- 42
        41716 => X"3D",  -- 61
        41717 => X"55",  -- 85
        41718 => X"73",  -- 115
        41719 => X"88",  -- 136
        41720 => X"96",  -- 150
        41721 => X"85",  -- 133
        41722 => X"7C",  -- 124
        41723 => X"77",  -- 119
        41724 => X"72",  -- 114
        41725 => X"71",  -- 113
        41726 => X"75",  -- 117
        41727 => X"72",  -- 114
        41728 => X"5D",  -- 93
        41729 => X"71",  -- 113
        41730 => X"7C",  -- 124
        41731 => X"7D",  -- 125
        41732 => X"87",  -- 135
        41733 => X"86",  -- 134
        41734 => X"75",  -- 117
        41735 => X"67",  -- 103
        41736 => X"52",  -- 82
        41737 => X"2D",  -- 45
        41738 => X"2E",  -- 46
        41739 => X"63",  -- 99
        41740 => X"B0",  -- 176
        41741 => X"D5",  -- 213
        41742 => X"CA",  -- 202
        41743 => X"C9",  -- 201
        41744 => X"D9",  -- 217
        41745 => X"A8",  -- 168
        41746 => X"63",  -- 99
        41747 => X"8E",  -- 142
        41748 => X"C7",  -- 199
        41749 => X"D1",  -- 209
        41750 => X"D2",  -- 210
        41751 => X"DC",  -- 220
        41752 => X"DE",  -- 222
        41753 => X"D5",  -- 213
        41754 => X"A6",  -- 166
        41755 => X"46",  -- 70
        41756 => X"1F",  -- 31
        41757 => X"28",  -- 40
        41758 => X"1E",  -- 30
        41759 => X"47",  -- 71
        41760 => X"79",  -- 121
        41761 => X"BD",  -- 189
        41762 => X"D2",  -- 210
        41763 => X"C3",  -- 195
        41764 => X"B7",  -- 183
        41765 => X"A6",  -- 166
        41766 => X"A6",  -- 166
        41767 => X"AD",  -- 173
        41768 => X"AF",  -- 175
        41769 => X"B0",  -- 176
        41770 => X"C1",  -- 193
        41771 => X"C4",  -- 196
        41772 => X"D8",  -- 216
        41773 => X"D2",  -- 210
        41774 => X"90",  -- 144
        41775 => X"71",  -- 113
        41776 => X"84",  -- 132
        41777 => X"82",  -- 130
        41778 => X"65",  -- 101
        41779 => X"6D",  -- 109
        41780 => X"70",  -- 112
        41781 => X"5F",  -- 95
        41782 => X"6A",  -- 106
        41783 => X"6A",  -- 106
        41784 => X"67",  -- 103
        41785 => X"5D",  -- 93
        41786 => X"52",  -- 82
        41787 => X"4E",  -- 78
        41788 => X"52",  -- 82
        41789 => X"57",  -- 87
        41790 => X"58",  -- 88
        41791 => X"56",  -- 86
        41792 => X"57",  -- 87
        41793 => X"5C",  -- 92
        41794 => X"5E",  -- 94
        41795 => X"5B",  -- 91
        41796 => X"59",  -- 89
        41797 => X"5C",  -- 92
        41798 => X"60",  -- 96
        41799 => X"62",  -- 98
        41800 => X"5F",  -- 95
        41801 => X"5D",  -- 93
        41802 => X"60",  -- 96
        41803 => X"64",  -- 100
        41804 => X"61",  -- 97
        41805 => X"59",  -- 89
        41806 => X"57",  -- 87
        41807 => X"5A",  -- 90
        41808 => X"61",  -- 97
        41809 => X"5F",  -- 95
        41810 => X"5B",  -- 91
        41811 => X"57",  -- 87
        41812 => X"57",  -- 87
        41813 => X"58",  -- 88
        41814 => X"56",  -- 86
        41815 => X"51",  -- 81
        41816 => X"47",  -- 71
        41817 => X"4B",  -- 75
        41818 => X"50",  -- 80
        41819 => X"51",  -- 81
        41820 => X"4F",  -- 79
        41821 => X"4A",  -- 74
        41822 => X"46",  -- 70
        41823 => X"44",  -- 68
        41824 => X"47",  -- 71
        41825 => X"4A",  -- 74
        41826 => X"44",  -- 68
        41827 => X"3F",  -- 63
        41828 => X"43",  -- 67
        41829 => X"43",  -- 67
        41830 => X"48",  -- 72
        41831 => X"52",  -- 82
        41832 => X"6D",  -- 109
        41833 => X"74",  -- 116
        41834 => X"7E",  -- 126
        41835 => X"87",  -- 135
        41836 => X"94",  -- 148
        41837 => X"A4",  -- 164
        41838 => X"B0",  -- 176
        41839 => X"B4",  -- 180
        41840 => X"BF",  -- 191
        41841 => X"BD",  -- 189
        41842 => X"C6",  -- 198
        41843 => X"C3",  -- 195
        41844 => X"C5",  -- 197
        41845 => X"CC",  -- 204
        41846 => X"BE",  -- 190
        41847 => X"BB",  -- 187
        41848 => X"C3",  -- 195
        41849 => X"BA",  -- 186
        41850 => X"B8",  -- 184
        41851 => X"B2",  -- 178
        41852 => X"A2",  -- 162
        41853 => X"A6",  -- 166
        41854 => X"AE",  -- 174
        41855 => X"A6",  -- 166
        41856 => X"A3",  -- 163
        41857 => X"9C",  -- 156
        41858 => X"A1",  -- 161
        41859 => X"AB",  -- 171
        41860 => X"A4",  -- 164
        41861 => X"9A",  -- 154
        41862 => X"9E",  -- 158
        41863 => X"A6",  -- 166
        41864 => X"9E",  -- 158
        41865 => X"9B",  -- 155
        41866 => X"97",  -- 151
        41867 => X"94",  -- 148
        41868 => X"95",  -- 149
        41869 => X"96",  -- 150
        41870 => X"9B",  -- 155
        41871 => X"9E",  -- 158
        41872 => X"A8",  -- 168
        41873 => X"B0",  -- 176
        41874 => X"B2",  -- 178
        41875 => X"AB",  -- 171
        41876 => X"A8",  -- 168
        41877 => X"AE",  -- 174
        41878 => X"B2",  -- 178
        41879 => X"B3",  -- 179
        41880 => X"AA",  -- 170
        41881 => X"AA",  -- 170
        41882 => X"AB",  -- 171
        41883 => X"AE",  -- 174
        41884 => X"B3",  -- 179
        41885 => X"B8",  -- 184
        41886 => X"BE",  -- 190
        41887 => X"C6",  -- 198
        41888 => X"C7",  -- 199
        41889 => X"CA",  -- 202
        41890 => X"CA",  -- 202
        41891 => X"C8",  -- 200
        41892 => X"C6",  -- 198
        41893 => X"C5",  -- 197
        41894 => X"BE",  -- 190
        41895 => X"B7",  -- 183
        41896 => X"A4",  -- 164
        41897 => X"99",  -- 153
        41898 => X"9A",  -- 154
        41899 => X"A4",  -- 164
        41900 => X"AC",  -- 172
        41901 => X"B3",  -- 179
        41902 => X"B0",  -- 176
        41903 => X"A4",  -- 164
        41904 => X"9F",  -- 159
        41905 => X"8B",  -- 139
        41906 => X"94",  -- 148
        41907 => X"8A",  -- 138
        41908 => X"7F",  -- 127
        41909 => X"78",  -- 120
        41910 => X"59",  -- 89
        41911 => X"52",  -- 82
        41912 => X"62",  -- 98
        41913 => X"76",  -- 118
        41914 => X"97",  -- 151
        41915 => X"A8",  -- 168
        41916 => X"9A",  -- 154
        41917 => X"77",  -- 119
        41918 => X"5A",  -- 90
        41919 => X"4F",  -- 79
        41920 => X"68",  -- 104
        41921 => X"64",  -- 100
        41922 => X"60",  -- 96
        41923 => X"62",  -- 98
        41924 => X"6D",  -- 109
        41925 => X"7C",  -- 124
        41926 => X"8A",  -- 138
        41927 => X"92",  -- 146
        41928 => X"96",  -- 150
        41929 => X"90",  -- 144
        41930 => X"87",  -- 135
        41931 => X"80",  -- 128
        41932 => X"79",  -- 121
        41933 => X"6F",  -- 111
        41934 => X"62",  -- 98
        41935 => X"59",  -- 89
        41936 => X"52",  -- 82
        41937 => X"50",  -- 80
        41938 => X"4C",  -- 76
        41939 => X"4B",  -- 75
        41940 => X"4C",  -- 76
        41941 => X"4E",  -- 78
        41942 => X"4F",  -- 79
        41943 => X"50",  -- 80
        41944 => X"52",  -- 82
        41945 => X"5A",  -- 90
        41946 => X"61",  -- 97
        41947 => X"63",  -- 99
        41948 => X"64",  -- 100
        41949 => X"65",  -- 101
        41950 => X"5A",  -- 90
        41951 => X"48",  -- 72
        41952 => X"55",  -- 85
        41953 => X"6A",  -- 106
        41954 => X"5D",  -- 93
        41955 => X"2C",  -- 44
        41956 => X"1A",  -- 26
        41957 => X"12",  -- 18
        41958 => X"18",  -- 24
        41959 => X"46",  -- 70
        41960 => X"88",  -- 136
        41961 => X"90",  -- 144
        41962 => X"93",  -- 147
        41963 => X"8D",  -- 141
        41964 => X"85",  -- 133
        41965 => X"47",  -- 71
        41966 => X"21",  -- 33
        41967 => X"66",  -- 102
        41968 => X"88",  -- 136
        41969 => X"91",  -- 145
        41970 => X"85",  -- 133
        41971 => X"5E",  -- 94
        41972 => X"1E",  -- 30
        41973 => X"16",  -- 22
        41974 => X"3A",  -- 58
        41975 => X"26",  -- 38
        41976 => X"2B",  -- 43
        41977 => X"52",  -- 82
        41978 => X"67",  -- 103
        41979 => X"5F",  -- 95
        41980 => X"5C",  -- 92
        41981 => X"60",  -- 96
        41982 => X"5D",  -- 93
        41983 => X"59",  -- 89
        41984 => X"5E",  -- 94
        41985 => X"5E",  -- 94
        41986 => X"5A",  -- 90
        41987 => X"65",  -- 101
        41988 => X"68",  -- 104
        41989 => X"67",  -- 103
        41990 => X"69",  -- 105
        41991 => X"4C",  -- 76
        41992 => X"31",  -- 49
        41993 => X"20",  -- 32
        41994 => X"13",  -- 19
        41995 => X"24",  -- 36
        41996 => X"3C",  -- 60
        41997 => X"3E",  -- 62
        41998 => X"30",  -- 48
        41999 => X"2E",  -- 46
        42000 => X"31",  -- 49
        42001 => X"2E",  -- 46
        42002 => X"2F",  -- 47
        42003 => X"34",  -- 52
        42004 => X"3A",  -- 58
        42005 => X"3E",  -- 62
        42006 => X"46",  -- 70
        42007 => X"4E",  -- 78
        42008 => X"45",  -- 69
        42009 => X"4A",  -- 74
        42010 => X"50",  -- 80
        42011 => X"51",  -- 81
        42012 => X"51",  -- 81
        42013 => X"51",  -- 81
        42014 => X"4F",  -- 79
        42015 => X"4D",  -- 77
        42016 => X"44",  -- 68
        42017 => X"57",  -- 87
        42018 => X"5C",  -- 92
        42019 => X"6C",  -- 108
        42020 => X"72",  -- 114
        42021 => X"7D",  -- 125
        42022 => X"6F",  -- 111
        42023 => X"6E",  -- 110
        42024 => X"6B",  -- 107
        42025 => X"6C",  -- 108
        42026 => X"68",  -- 104
        42027 => X"5F",  -- 95
        42028 => X"5C",  -- 92
        42029 => X"5F",  -- 95
        42030 => X"60",  -- 96
        42031 => X"5D",  -- 93
        42032 => X"4F",  -- 79
        42033 => X"2C",  -- 44
        42034 => X"29",  -- 41
        42035 => X"2A",  -- 42
        42036 => X"36",  -- 54
        42037 => X"55",  -- 85
        42038 => X"6C",  -- 108
        42039 => X"8A",  -- 138
        42040 => X"95",  -- 149
        42041 => X"86",  -- 134
        42042 => X"7C",  -- 124
        42043 => X"78",  -- 120
        42044 => X"72",  -- 114
        42045 => X"7A",  -- 122
        42046 => X"85",  -- 133
        42047 => X"86",  -- 134
        42048 => X"59",  -- 89
        42049 => X"65",  -- 101
        42050 => X"71",  -- 113
        42051 => X"78",  -- 120
        42052 => X"82",  -- 130
        42053 => X"6D",  -- 109
        42054 => X"39",  -- 57
        42055 => X"1F",  -- 31
        42056 => X"1E",  -- 30
        42057 => X"5A",  -- 90
        42058 => X"95",  -- 149
        42059 => X"B6",  -- 182
        42060 => X"CF",  -- 207
        42061 => X"D6",  -- 214
        42062 => X"CD",  -- 205
        42063 => X"D5",  -- 213
        42064 => X"D7",  -- 215
        42065 => X"89",  -- 137
        42066 => X"67",  -- 103
        42067 => X"A4",  -- 164
        42068 => X"D2",  -- 210
        42069 => X"CF",  -- 207
        42070 => X"D0",  -- 208
        42071 => X"DE",  -- 222
        42072 => X"E0",  -- 224
        42073 => X"DF",  -- 223
        42074 => X"C4",  -- 196
        42075 => X"62",  -- 98
        42076 => X"16",  -- 22
        42077 => X"1D",  -- 29
        42078 => X"19",  -- 25
        42079 => X"46",  -- 70
        42080 => X"6E",  -- 110
        42081 => X"AF",  -- 175
        42082 => X"CB",  -- 203
        42083 => X"C5",  -- 197
        42084 => X"BB",  -- 187
        42085 => X"AF",  -- 175
        42086 => X"A8",  -- 168
        42087 => X"9A",  -- 154
        42088 => X"B7",  -- 183
        42089 => X"BE",  -- 190
        42090 => X"C3",  -- 195
        42091 => X"C0",  -- 192
        42092 => X"CD",  -- 205
        42093 => X"D5",  -- 213
        42094 => X"AE",  -- 174
        42095 => X"7C",  -- 124
        42096 => X"7A",  -- 122
        42097 => X"7E",  -- 126
        42098 => X"65",  -- 101
        42099 => X"61",  -- 97
        42100 => X"66",  -- 102
        42101 => X"5A",  -- 90
        42102 => X"5F",  -- 95
        42103 => X"65",  -- 101
        42104 => X"67",  -- 103
        42105 => X"5E",  -- 94
        42106 => X"55",  -- 85
        42107 => X"54",  -- 84
        42108 => X"59",  -- 89
        42109 => X"5C",  -- 92
        42110 => X"59",  -- 89
        42111 => X"55",  -- 85
        42112 => X"56",  -- 86
        42113 => X"5B",  -- 91
        42114 => X"5F",  -- 95
        42115 => X"5D",  -- 93
        42116 => X"59",  -- 89
        42117 => X"57",  -- 87
        42118 => X"59",  -- 89
        42119 => X"5B",  -- 91
        42120 => X"5A",  -- 90
        42121 => X"57",  -- 87
        42122 => X"59",  -- 89
        42123 => X"5F",  -- 95
        42124 => X"61",  -- 97
        42125 => X"5C",  -- 92
        42126 => X"58",  -- 88
        42127 => X"57",  -- 87
        42128 => X"5F",  -- 95
        42129 => X"5C",  -- 92
        42130 => X"58",  -- 88
        42131 => X"55",  -- 85
        42132 => X"54",  -- 84
        42133 => X"54",  -- 84
        42134 => X"52",  -- 82
        42135 => X"50",  -- 80
        42136 => X"45",  -- 69
        42137 => X"49",  -- 73
        42138 => X"4C",  -- 76
        42139 => X"4D",  -- 77
        42140 => X"4B",  -- 75
        42141 => X"47",  -- 71
        42142 => X"44",  -- 68
        42143 => X"44",  -- 68
        42144 => X"44",  -- 68
        42145 => X"46",  -- 70
        42146 => X"41",  -- 65
        42147 => X"3E",  -- 62
        42148 => X"42",  -- 66
        42149 => X"43",  -- 67
        42150 => X"4A",  -- 74
        42151 => X"57",  -- 87
        42152 => X"73",  -- 115
        42153 => X"79",  -- 121
        42154 => X"82",  -- 130
        42155 => X"8C",  -- 140
        42156 => X"99",  -- 153
        42157 => X"A8",  -- 168
        42158 => X"AF",  -- 175
        42159 => X"AE",  -- 174
        42160 => X"B6",  -- 182
        42161 => X"B6",  -- 182
        42162 => X"BD",  -- 189
        42163 => X"B9",  -- 185
        42164 => X"BD",  -- 189
        42165 => X"C7",  -- 199
        42166 => X"BF",  -- 191
        42167 => X"BC",  -- 188
        42168 => X"BD",  -- 189
        42169 => X"B2",  -- 178
        42170 => X"B8",  -- 184
        42171 => X"B3",  -- 179
        42172 => X"A1",  -- 161
        42173 => X"AB",  -- 171
        42174 => X"B6",  -- 182
        42175 => X"A7",  -- 167
        42176 => X"B2",  -- 178
        42177 => X"A1",  -- 161
        42178 => X"A8",  -- 168
        42179 => X"AE",  -- 174
        42180 => X"9E",  -- 158
        42181 => X"95",  -- 149
        42182 => X"9D",  -- 157
        42183 => X"A2",  -- 162
        42184 => X"9A",  -- 154
        42185 => X"95",  -- 149
        42186 => X"92",  -- 146
        42187 => X"93",  -- 147
        42188 => X"98",  -- 152
        42189 => X"9E",  -- 158
        42190 => X"A3",  -- 163
        42191 => X"A5",  -- 165
        42192 => X"A7",  -- 167
        42193 => X"AD",  -- 173
        42194 => X"AD",  -- 173
        42195 => X"A7",  -- 167
        42196 => X"A6",  -- 166
        42197 => X"AE",  -- 174
        42198 => X"B4",  -- 180
        42199 => X"B4",  -- 180
        42200 => X"AE",  -- 174
        42201 => X"AB",  -- 171
        42202 => X"A7",  -- 167
        42203 => X"AB",  -- 171
        42204 => X"B5",  -- 181
        42205 => X"BC",  -- 188
        42206 => X"C3",  -- 195
        42207 => X"C6",  -- 198
        42208 => X"C4",  -- 196
        42209 => X"CA",  -- 202
        42210 => X"CC",  -- 204
        42211 => X"CB",  -- 203
        42212 => X"C9",  -- 201
        42213 => X"C7",  -- 199
        42214 => X"C2",  -- 194
        42215 => X"BC",  -- 188
        42216 => X"AE",  -- 174
        42217 => X"9F",  -- 159
        42218 => X"9B",  -- 155
        42219 => X"A0",  -- 160
        42220 => X"A6",  -- 166
        42221 => X"AE",  -- 174
        42222 => X"AD",  -- 173
        42223 => X"A2",  -- 162
        42224 => X"9D",  -- 157
        42225 => X"83",  -- 131
        42226 => X"72",  -- 114
        42227 => X"86",  -- 134
        42228 => X"75",  -- 117
        42229 => X"62",  -- 98
        42230 => X"6D",  -- 109
        42231 => X"54",  -- 84
        42232 => X"62",  -- 98
        42233 => X"6B",  -- 107
        42234 => X"82",  -- 130
        42235 => X"99",  -- 153
        42236 => X"A0",  -- 160
        42237 => X"8B",  -- 139
        42238 => X"69",  -- 105
        42239 => X"53",  -- 83
        42240 => X"6C",  -- 108
        42241 => X"69",  -- 105
        42242 => X"66",  -- 102
        42243 => X"65",  -- 101
        42244 => X"6B",  -- 107
        42245 => X"78",  -- 120
        42246 => X"89",  -- 137
        42247 => X"95",  -- 149
        42248 => X"9A",  -- 154
        42249 => X"96",  -- 150
        42250 => X"91",  -- 145
        42251 => X"8A",  -- 138
        42252 => X"81",  -- 129
        42253 => X"75",  -- 117
        42254 => X"69",  -- 105
        42255 => X"60",  -- 96
        42256 => X"58",  -- 88
        42257 => X"54",  -- 84
        42258 => X"4F",  -- 79
        42259 => X"4E",  -- 78
        42260 => X"4F",  -- 79
        42261 => X"50",  -- 80
        42262 => X"51",  -- 81
        42263 => X"50",  -- 80
        42264 => X"52",  -- 82
        42265 => X"5F",  -- 95
        42266 => X"66",  -- 102
        42267 => X"65",  -- 101
        42268 => X"63",  -- 99
        42269 => X"5C",  -- 92
        42270 => X"50",  -- 80
        42271 => X"45",  -- 69
        42272 => X"5D",  -- 93
        42273 => X"71",  -- 113
        42274 => X"63",  -- 99
        42275 => X"39",  -- 57
        42276 => X"26",  -- 38
        42277 => X"1A",  -- 26
        42278 => X"18",  -- 24
        42279 => X"43",  -- 67
        42280 => X"82",  -- 130
        42281 => X"83",  -- 131
        42282 => X"95",  -- 149
        42283 => X"8A",  -- 138
        42284 => X"6E",  -- 110
        42285 => X"43",  -- 67
        42286 => X"23",  -- 35
        42287 => X"43",  -- 67
        42288 => X"87",  -- 135
        42289 => X"93",  -- 147
        42290 => X"8B",  -- 139
        42291 => X"86",  -- 134
        42292 => X"5E",  -- 94
        42293 => X"2E",  -- 46
        42294 => X"3E",  -- 62
        42295 => X"54",  -- 84
        42296 => X"5D",  -- 93
        42297 => X"65",  -- 101
        42298 => X"6B",  -- 107
        42299 => X"6C",  -- 108
        42300 => X"61",  -- 97
        42301 => X"4C",  -- 76
        42302 => X"4E",  -- 78
        42303 => X"63",  -- 99
        42304 => X"63",  -- 99
        42305 => X"5D",  -- 93
        42306 => X"59",  -- 89
        42307 => X"64",  -- 100
        42308 => X"6A",  -- 106
        42309 => X"67",  -- 103
        42310 => X"5D",  -- 93
        42311 => X"46",  -- 70
        42312 => X"30",  -- 48
        42313 => X"21",  -- 33
        42314 => X"14",  -- 20
        42315 => X"21",  -- 33
        42316 => X"34",  -- 52
        42317 => X"32",  -- 50
        42318 => X"29",  -- 41
        42319 => X"2C",  -- 44
        42320 => X"31",  -- 49
        42321 => X"30",  -- 48
        42322 => X"31",  -- 49
        42323 => X"34",  -- 52
        42324 => X"39",  -- 57
        42325 => X"3D",  -- 61
        42326 => X"47",  -- 71
        42327 => X"4E",  -- 78
        42328 => X"57",  -- 87
        42329 => X"4F",  -- 79
        42330 => X"4D",  -- 77
        42331 => X"50",  -- 80
        42332 => X"4F",  -- 79
        42333 => X"4B",  -- 75
        42334 => X"4D",  -- 77
        42335 => X"56",  -- 86
        42336 => X"4F",  -- 79
        42337 => X"5E",  -- 94
        42338 => X"63",  -- 99
        42339 => X"77",  -- 119
        42340 => X"72",  -- 114
        42341 => X"6E",  -- 110
        42342 => X"5F",  -- 95
        42343 => X"69",  -- 105
        42344 => X"66",  -- 102
        42345 => X"6C",  -- 108
        42346 => X"6B",  -- 107
        42347 => X"61",  -- 97
        42348 => X"5E",  -- 94
        42349 => X"62",  -- 98
        42350 => X"60",  -- 96
        42351 => X"59",  -- 89
        42352 => X"41",  -- 65
        42353 => X"27",  -- 39
        42354 => X"30",  -- 48
        42355 => X"30",  -- 48
        42356 => X"3A",  -- 58
        42357 => X"57",  -- 87
        42358 => X"65",  -- 101
        42359 => X"7F",  -- 127
        42360 => X"91",  -- 145
        42361 => X"88",  -- 136
        42362 => X"82",  -- 130
        42363 => X"7C",  -- 124
        42364 => X"78",  -- 120
        42365 => X"82",  -- 130
        42366 => X"8E",  -- 142
        42367 => X"8E",  -- 142
        42368 => X"83",  -- 131
        42369 => X"7B",  -- 123
        42370 => X"75",  -- 117
        42371 => X"6C",  -- 108
        42372 => X"68",  -- 104
        42373 => X"47",  -- 71
        42374 => X"16",  -- 22
        42375 => X"15",  -- 21
        42376 => X"39",  -- 57
        42377 => X"8D",  -- 141
        42378 => X"C5",  -- 197
        42379 => X"D1",  -- 209
        42380 => X"D0",  -- 208
        42381 => X"CE",  -- 206
        42382 => X"CD",  -- 205
        42383 => X"CD",  -- 205
        42384 => X"BA",  -- 186
        42385 => X"62",  -- 98
        42386 => X"61",  -- 97
        42387 => X"A6",  -- 166
        42388 => X"CE",  -- 206
        42389 => X"C8",  -- 200
        42390 => X"C8",  -- 200
        42391 => X"D1",  -- 209
        42392 => X"D5",  -- 213
        42393 => X"DB",  -- 219
        42394 => X"DA",  -- 218
        42395 => X"96",  -- 150
        42396 => X"30",  -- 48
        42397 => X"1E",  -- 30
        42398 => X"12",  -- 18
        42399 => X"34",  -- 52
        42400 => X"6B",  -- 107
        42401 => X"A1",  -- 161
        42402 => X"C7",  -- 199
        42403 => X"C9",  -- 201
        42404 => X"B4",  -- 180
        42405 => X"B3",  -- 179
        42406 => X"AF",  -- 175
        42407 => X"86",  -- 134
        42408 => X"AA",  -- 170
        42409 => X"C7",  -- 199
        42410 => X"BF",  -- 191
        42411 => X"C1",  -- 193
        42412 => X"BD",  -- 189
        42413 => X"BC",  -- 188
        42414 => X"BE",  -- 190
        42415 => X"89",  -- 137
        42416 => X"71",  -- 113
        42417 => X"77",  -- 119
        42418 => X"73",  -- 115
        42419 => X"5C",  -- 92
        42420 => X"60",  -- 96
        42421 => X"65",  -- 101
        42422 => X"55",  -- 85
        42423 => X"5A",  -- 90
        42424 => X"60",  -- 96
        42425 => X"5A",  -- 90
        42426 => X"54",  -- 84
        42427 => X"55",  -- 85
        42428 => X"5A",  -- 90
        42429 => X"5D",  -- 93
        42430 => X"5A",  -- 90
        42431 => X"56",  -- 86
        42432 => X"55",  -- 85
        42433 => X"59",  -- 89
        42434 => X"5D",  -- 93
        42435 => X"5E",  -- 94
        42436 => X"59",  -- 89
        42437 => X"54",  -- 84
        42438 => X"52",  -- 82
        42439 => X"53",  -- 83
        42440 => X"57",  -- 87
        42441 => X"54",  -- 84
        42442 => X"53",  -- 83
        42443 => X"58",  -- 88
        42444 => X"5D",  -- 93
        42445 => X"5D",  -- 93
        42446 => X"5A",  -- 90
        42447 => X"59",  -- 89
        42448 => X"5C",  -- 92
        42449 => X"5A",  -- 90
        42450 => X"57",  -- 87
        42451 => X"55",  -- 85
        42452 => X"53",  -- 83
        42453 => X"51",  -- 81
        42454 => X"50",  -- 80
        42455 => X"50",  -- 80
        42456 => X"47",  -- 71
        42457 => X"48",  -- 72
        42458 => X"49",  -- 73
        42459 => X"49",  -- 73
        42460 => X"47",  -- 71
        42461 => X"45",  -- 69
        42462 => X"44",  -- 68
        42463 => X"45",  -- 69
        42464 => X"42",  -- 66
        42465 => X"43",  -- 67
        42466 => X"3F",  -- 63
        42467 => X"3D",  -- 61
        42468 => X"42",  -- 66
        42469 => X"42",  -- 66
        42470 => X"4B",  -- 75
        42471 => X"5B",  -- 91
        42472 => X"74",  -- 116
        42473 => X"7D",  -- 125
        42474 => X"87",  -- 135
        42475 => X"92",  -- 146
        42476 => X"A0",  -- 160
        42477 => X"AD",  -- 173
        42478 => X"B0",  -- 176
        42479 => X"AF",  -- 175
        42480 => X"AF",  -- 175
        42481 => X"B2",  -- 178
        42482 => X"BA",  -- 186
        42483 => X"B0",  -- 176
        42484 => X"B1",  -- 177
        42485 => X"BC",  -- 188
        42486 => X"B9",  -- 185
        42487 => X"BC",  -- 188
        42488 => X"BC",  -- 188
        42489 => X"B4",  -- 180
        42490 => X"BB",  -- 187
        42491 => X"B8",  -- 184
        42492 => X"A7",  -- 167
        42493 => X"AF",  -- 175
        42494 => X"B7",  -- 183
        42495 => X"A4",  -- 164
        42496 => X"B5",  -- 181
        42497 => X"A6",  -- 166
        42498 => X"A8",  -- 168
        42499 => X"AB",  -- 171
        42500 => X"9B",  -- 155
        42501 => X"97",  -- 151
        42502 => X"9F",  -- 159
        42503 => X"A0",  -- 160
        42504 => X"9F",  -- 159
        42505 => X"98",  -- 152
        42506 => X"94",  -- 148
        42507 => X"97",  -- 151
        42508 => X"A0",  -- 160
        42509 => X"A9",  -- 169
        42510 => X"AB",  -- 171
        42511 => X"AA",  -- 170
        42512 => X"AD",  -- 173
        42513 => X"AD",  -- 173
        42514 => X"A9",  -- 169
        42515 => X"A3",  -- 163
        42516 => X"A4",  -- 164
        42517 => X"AD",  -- 173
        42518 => X"B3",  -- 179
        42519 => X"B1",  -- 177
        42520 => X"B5",  -- 181
        42521 => X"AD",  -- 173
        42522 => X"A5",  -- 165
        42523 => X"A6",  -- 166
        42524 => X"B3",  -- 179
        42525 => X"C0",  -- 192
        42526 => X"C5",  -- 197
        42527 => X"C5",  -- 197
        42528 => X"C3",  -- 195
        42529 => X"CA",  -- 202
        42530 => X"CE",  -- 206
        42531 => X"CD",  -- 205
        42532 => X"CA",  -- 202
        42533 => X"C5",  -- 197
        42534 => X"BD",  -- 189
        42535 => X"B6",  -- 182
        42536 => X"B2",  -- 178
        42537 => X"A5",  -- 165
        42538 => X"A1",  -- 161
        42539 => X"A3",  -- 163
        42540 => X"A2",  -- 162
        42541 => X"A6",  -- 166
        42542 => X"A5",  -- 165
        42543 => X"9C",  -- 156
        42544 => X"8B",  -- 139
        42545 => X"90",  -- 144
        42546 => X"63",  -- 99
        42547 => X"5C",  -- 92
        42548 => X"68",  -- 104
        42549 => X"5A",  -- 90
        42550 => X"61",  -- 97
        42551 => X"67",  -- 103
        42552 => X"6B",  -- 107
        42553 => X"6E",  -- 110
        42554 => X"76",  -- 118
        42555 => X"7E",  -- 126
        42556 => X"89",  -- 137
        42557 => X"88",  -- 136
        42558 => X"77",  -- 119
        42559 => X"64",  -- 100
        42560 => X"6B",  -- 107
        42561 => X"6C",  -- 108
        42562 => X"6C",  -- 108
        42563 => X"6B",  -- 107
        42564 => X"6B",  -- 107
        42565 => X"73",  -- 115
        42566 => X"80",  -- 128
        42567 => X"8A",  -- 138
        42568 => X"8D",  -- 141
        42569 => X"8E",  -- 142
        42570 => X"8E",  -- 142
        42571 => X"89",  -- 137
        42572 => X"80",  -- 128
        42573 => X"75",  -- 117
        42574 => X"6C",  -- 108
        42575 => X"65",  -- 101
        42576 => X"5D",  -- 93
        42577 => X"59",  -- 89
        42578 => X"55",  -- 85
        42579 => X"52",  -- 82
        42580 => X"52",  -- 82
        42581 => X"52",  -- 82
        42582 => X"51",  -- 81
        42583 => X"50",  -- 80
        42584 => X"51",  -- 81
        42585 => X"61",  -- 97
        42586 => X"68",  -- 104
        42587 => X"62",  -- 98
        42588 => X"5D",  -- 93
        42589 => X"52",  -- 82
        42590 => X"46",  -- 70
        42591 => X"47",  -- 71
        42592 => X"69",  -- 105
        42593 => X"71",  -- 113
        42594 => X"66",  -- 102
        42595 => X"45",  -- 69
        42596 => X"31",  -- 49
        42597 => X"21",  -- 33
        42598 => X"1B",  -- 27
        42599 => X"3D",  -- 61
        42600 => X"7A",  -- 122
        42601 => X"7D",  -- 125
        42602 => X"8E",  -- 142
        42603 => X"81",  -- 129
        42604 => X"54",  -- 84
        42605 => X"2E",  -- 46
        42606 => X"1A",  -- 26
        42607 => X"18",  -- 24
        42608 => X"5C",  -- 92
        42609 => X"8D",  -- 141
        42610 => X"96",  -- 150
        42611 => X"91",  -- 145
        42612 => X"8E",  -- 142
        42613 => X"75",  -- 117
        42614 => X"66",  -- 102
        42615 => X"69",  -- 105
        42616 => X"44",  -- 68
        42617 => X"4B",  -- 75
        42618 => X"4F",  -- 79
        42619 => X"55",  -- 85
        42620 => X"54",  -- 84
        42621 => X"4C",  -- 76
        42622 => X"51",  -- 81
        42623 => X"61",  -- 97
        42624 => X"62",  -- 98
        42625 => X"62",  -- 98
        42626 => X"61",  -- 97
        42627 => X"65",  -- 101
        42628 => X"66",  -- 102
        42629 => X"5B",  -- 91
        42630 => X"4C",  -- 76
        42631 => X"40",  -- 64
        42632 => X"2D",  -- 45
        42633 => X"22",  -- 34
        42634 => X"15",  -- 21
        42635 => X"1A",  -- 26
        42636 => X"28",  -- 40
        42637 => X"28",  -- 40
        42638 => X"28",  -- 40
        42639 => X"31",  -- 49
        42640 => X"32",  -- 50
        42641 => X"30",  -- 48
        42642 => X"32",  -- 50
        42643 => X"36",  -- 54
        42644 => X"3A",  -- 58
        42645 => X"3F",  -- 63
        42646 => X"48",  -- 72
        42647 => X"50",  -- 80
        42648 => X"63",  -- 99
        42649 => X"57",  -- 87
        42650 => X"55",  -- 85
        42651 => X"5A",  -- 90
        42652 => X"54",  -- 84
        42653 => X"44",  -- 68
        42654 => X"40",  -- 64
        42655 => X"47",  -- 71
        42656 => X"60",  -- 96
        42657 => X"67",  -- 103
        42658 => X"68",  -- 104
        42659 => X"7D",  -- 125
        42660 => X"77",  -- 119
        42661 => X"72",  -- 114
        42662 => X"68",  -- 104
        42663 => X"7A",  -- 122
        42664 => X"66",  -- 102
        42665 => X"6A",  -- 106
        42666 => X"69",  -- 105
        42667 => X"61",  -- 97
        42668 => X"5C",  -- 92
        42669 => X"5C",  -- 92
        42670 => X"57",  -- 87
        42671 => X"4D",  -- 77
        42672 => X"42",  -- 66
        42673 => X"27",  -- 39
        42674 => X"2A",  -- 42
        42675 => X"2C",  -- 44
        42676 => X"3A",  -- 58
        42677 => X"59",  -- 89
        42678 => X"65",  -- 101
        42679 => X"75",  -- 117
        42680 => X"8A",  -- 138
        42681 => X"88",  -- 136
        42682 => X"89",  -- 137
        42683 => X"85",  -- 133
        42684 => X"7E",  -- 126
        42685 => X"83",  -- 131
        42686 => X"88",  -- 136
        42687 => X"84",  -- 132
        42688 => X"8A",  -- 138
        42689 => X"83",  -- 131
        42690 => X"84",  -- 132
        42691 => X"73",  -- 115
        42692 => X"67",  -- 103
        42693 => X"40",  -- 64
        42694 => X"12",  -- 18
        42695 => X"2A",  -- 42
        42696 => X"6E",  -- 110
        42697 => X"A4",  -- 164
        42698 => X"C8",  -- 200
        42699 => X"D2",  -- 210
        42700 => X"CF",  -- 207
        42701 => X"C6",  -- 198
        42702 => X"CC",  -- 204
        42703 => X"CA",  -- 202
        42704 => X"9B",  -- 155
        42705 => X"4D",  -- 77
        42706 => X"6B",  -- 107
        42707 => X"A6",  -- 166
        42708 => X"C8",  -- 200
        42709 => X"CB",  -- 203
        42710 => X"C7",  -- 199
        42711 => X"CA",  -- 202
        42712 => X"D3",  -- 211
        42713 => X"CF",  -- 207
        42714 => X"CF",  -- 207
        42715 => X"AD",  -- 173
        42716 => X"42",  -- 66
        42717 => X"21",  -- 33
        42718 => X"1B",  -- 27
        42719 => X"2B",  -- 43
        42720 => X"6B",  -- 107
        42721 => X"98",  -- 152
        42722 => X"C0",  -- 192
        42723 => X"C5",  -- 197
        42724 => X"AA",  -- 170
        42725 => X"AD",  -- 173
        42726 => X"B5",  -- 181
        42727 => X"8F",  -- 143
        42728 => X"9C",  -- 156
        42729 => X"C6",  -- 198
        42730 => X"BF",  -- 191
        42731 => X"CB",  -- 203
        42732 => X"BA",  -- 186
        42733 => X"A5",  -- 165
        42734 => X"B5",  -- 181
        42735 => X"89",  -- 137
        42736 => X"6B",  -- 107
        42737 => X"6E",  -- 110
        42738 => X"79",  -- 121
        42739 => X"5F",  -- 95
        42740 => X"5F",  -- 95
        42741 => X"6E",  -- 110
        42742 => X"56",  -- 86
        42743 => X"53",  -- 83
        42744 => X"5A",  -- 90
        42745 => X"54",  -- 84
        42746 => X"50",  -- 80
        42747 => X"4F",  -- 79
        42748 => X"53",  -- 83
        42749 => X"59",  -- 89
        42750 => X"5B",  -- 91
        42751 => X"5C",  -- 92
        42752 => X"57",  -- 87
        42753 => X"57",  -- 87
        42754 => X"59",  -- 89
        42755 => X"5B",  -- 91
        42756 => X"58",  -- 88
        42757 => X"52",  -- 82
        42758 => X"4F",  -- 79
        42759 => X"4F",  -- 79
        42760 => X"56",  -- 86
        42761 => X"52",  -- 82
        42762 => X"50",  -- 80
        42763 => X"52",  -- 82
        42764 => X"57",  -- 87
        42765 => X"5A",  -- 90
        42766 => X"5A",  -- 90
        42767 => X"58",  -- 88
        42768 => X"59",  -- 89
        42769 => X"56",  -- 86
        42770 => X"55",  -- 85
        42771 => X"55",  -- 85
        42772 => X"53",  -- 83
        42773 => X"50",  -- 80
        42774 => X"4E",  -- 78
        42775 => X"4F",  -- 79
        42776 => X"47",  -- 71
        42777 => X"48",  -- 72
        42778 => X"48",  -- 72
        42779 => X"46",  -- 70
        42780 => X"44",  -- 68
        42781 => X"42",  -- 66
        42782 => X"42",  -- 66
        42783 => X"44",  -- 68
        42784 => X"42",  -- 66
        42785 => X"41",  -- 65
        42786 => X"3E",  -- 62
        42787 => X"3D",  -- 61
        42788 => X"42",  -- 66
        42789 => X"42",  -- 66
        42790 => X"4D",  -- 77
        42791 => X"60",  -- 96
        42792 => X"74",  -- 116
        42793 => X"7F",  -- 127
        42794 => X"8B",  -- 139
        42795 => X"9A",  -- 154
        42796 => X"A7",  -- 167
        42797 => X"B1",  -- 177
        42798 => X"B5",  -- 181
        42799 => X"B1",  -- 177
        42800 => X"AC",  -- 172
        42801 => X"B2",  -- 178
        42802 => X"BB",  -- 187
        42803 => X"AA",  -- 170
        42804 => X"A5",  -- 165
        42805 => X"B1",  -- 177
        42806 => X"B3",  -- 179
        42807 => X"B8",  -- 184
        42808 => X"B8",  -- 184
        42809 => X"B1",  -- 177
        42810 => X"B7",  -- 183
        42811 => X"B8",  -- 184
        42812 => X"AF",  -- 175
        42813 => X"B3",  -- 179
        42814 => X"B6",  -- 182
        42815 => X"AA",  -- 170
        42816 => X"B3",  -- 179
        42817 => X"AD",  -- 173
        42818 => X"AB",  -- 171
        42819 => X"A9",  -- 169
        42820 => X"A2",  -- 162
        42821 => X"A1",  -- 161
        42822 => X"A6",  -- 166
        42823 => X"A5",  -- 165
        42824 => X"A6",  -- 166
        42825 => X"A0",  -- 160
        42826 => X"9C",  -- 156
        42827 => X"9E",  -- 158
        42828 => X"A3",  -- 163
        42829 => X"A8",  -- 168
        42830 => X"A8",  -- 168
        42831 => X"A5",  -- 165
        42832 => X"B2",  -- 178
        42833 => X"B2",  -- 178
        42834 => X"AB",  -- 171
        42835 => X"A3",  -- 163
        42836 => X"A5",  -- 165
        42837 => X"AE",  -- 174
        42838 => X"B1",  -- 177
        42839 => X"AC",  -- 172
        42840 => X"B6",  -- 182
        42841 => X"AF",  -- 175
        42842 => X"A8",  -- 168
        42843 => X"A6",  -- 166
        42844 => X"B1",  -- 177
        42845 => X"BE",  -- 190
        42846 => X"C4",  -- 196
        42847 => X"C6",  -- 198
        42848 => X"C4",  -- 196
        42849 => X"CA",  -- 202
        42850 => X"CE",  -- 206
        42851 => X"CD",  -- 205
        42852 => X"CA",  -- 202
        42853 => X"C4",  -- 196
        42854 => X"B8",  -- 184
        42855 => X"AD",  -- 173
        42856 => X"AF",  -- 175
        42857 => X"A6",  -- 166
        42858 => X"A5",  -- 165
        42859 => X"A5",  -- 165
        42860 => X"9F",  -- 159
        42861 => X"9F",  -- 159
        42862 => X"9D",  -- 157
        42863 => X"95",  -- 149
        42864 => X"8A",  -- 138
        42865 => X"80",  -- 128
        42866 => X"73",  -- 115
        42867 => X"4A",  -- 74
        42868 => X"46",  -- 70
        42869 => X"61",  -- 97
        42870 => X"62",  -- 98
        42871 => X"6F",  -- 111
        42872 => X"64",  -- 100
        42873 => X"71",  -- 113
        42874 => X"7D",  -- 125
        42875 => X"7C",  -- 124
        42876 => X"79",  -- 121
        42877 => X"75",  -- 117
        42878 => X"6C",  -- 108
        42879 => X"63",  -- 99
        42880 => X"66",  -- 102
        42881 => X"69",  -- 105
        42882 => X"6F",  -- 111
        42883 => X"70",  -- 112
        42884 => X"70",  -- 112
        42885 => X"72",  -- 114
        42886 => X"74",  -- 116
        42887 => X"76",  -- 118
        42888 => X"77",  -- 119
        42889 => X"7C",  -- 124
        42890 => X"80",  -- 128
        42891 => X"80",  -- 128
        42892 => X"7A",  -- 122
        42893 => X"72",  -- 114
        42894 => X"6B",  -- 107
        42895 => X"69",  -- 105
        42896 => X"60",  -- 96
        42897 => X"5C",  -- 92
        42898 => X"58",  -- 88
        42899 => X"57",  -- 87
        42900 => X"57",  -- 87
        42901 => X"56",  -- 86
        42902 => X"53",  -- 83
        42903 => X"4F",  -- 79
        42904 => X"4F",  -- 79
        42905 => X"5E",  -- 94
        42906 => X"60",  -- 96
        42907 => X"5D",  -- 93
        42908 => X"5A",  -- 90
        42909 => X"4E",  -- 78
        42910 => X"48",  -- 72
        42911 => X"57",  -- 87
        42912 => X"7B",  -- 123
        42913 => X"71",  -- 113
        42914 => X"65",  -- 101
        42915 => X"4D",  -- 77
        42916 => X"36",  -- 54
        42917 => X"22",  -- 34
        42918 => X"19",  -- 25
        42919 => X"33",  -- 51
        42920 => X"74",  -- 116
        42921 => X"7C",  -- 124
        42922 => X"7D",  -- 125
        42923 => X"71",  -- 113
        42924 => X"4A",  -- 74
        42925 => X"26",  -- 38
        42926 => X"20",  -- 32
        42927 => X"17",  -- 23
        42928 => X"29",  -- 41
        42929 => X"70",  -- 112
        42930 => X"94",  -- 148
        42931 => X"86",  -- 134
        42932 => X"8D",  -- 141
        42933 => X"92",  -- 146
        42934 => X"6C",  -- 108
        42935 => X"55",  -- 85
        42936 => X"20",  -- 32
        42937 => X"27",  -- 39
        42938 => X"25",  -- 37
        42939 => X"26",  -- 38
        42940 => X"39",  -- 57
        42941 => X"4B",  -- 75
        42942 => X"50",  -- 80
        42943 => X"54",  -- 84
        42944 => X"61",  -- 97
        42945 => X"62",  -- 98
        42946 => X"64",  -- 100
        42947 => X"60",  -- 96
        42948 => X"5F",  -- 95
        42949 => X"58",  -- 88
        42950 => X"44",  -- 68
        42951 => X"3D",  -- 61
        42952 => X"26",  -- 38
        42953 => X"21",  -- 33
        42954 => X"1A",  -- 26
        42955 => X"1E",  -- 30
        42956 => X"2C",  -- 44
        42957 => X"2E",  -- 46
        42958 => X"2D",  -- 45
        42959 => X"34",  -- 52
        42960 => X"32",  -- 50
        42961 => X"31",  -- 49
        42962 => X"34",  -- 52
        42963 => X"39",  -- 57
        42964 => X"3E",  -- 62
        42965 => X"42",  -- 66
        42966 => X"4B",  -- 75
        42967 => X"53",  -- 83
        42968 => X"4E",  -- 78
        42969 => X"4F",  -- 79
        42970 => X"56",  -- 86
        42971 => X"5F",  -- 95
        42972 => X"60",  -- 96
        42973 => X"58",  -- 88
        42974 => X"50",  -- 80
        42975 => X"4F",  -- 79
        42976 => X"61",  -- 97
        42977 => X"6B",  -- 107
        42978 => X"6D",  -- 109
        42979 => X"80",  -- 128
        42980 => X"80",  -- 128
        42981 => X"84",  -- 132
        42982 => X"7E",  -- 126
        42983 => X"8A",  -- 138
        42984 => X"70",  -- 112
        42985 => X"72",  -- 114
        42986 => X"6D",  -- 109
        42987 => X"65",  -- 101
        42988 => X"60",  -- 96
        42989 => X"5E",  -- 94
        42990 => X"5A",  -- 90
        42991 => X"54",  -- 84
        42992 => X"52",  -- 82
        42993 => X"3B",  -- 59
        42994 => X"34",  -- 52
        42995 => X"32",  -- 50
        42996 => X"3E",  -- 62
        42997 => X"5A",  -- 90
        42998 => X"6E",  -- 110
        42999 => X"7A",  -- 122
        43000 => X"81",  -- 129
        43001 => X"80",  -- 128
        43002 => X"84",  -- 132
        43003 => X"81",  -- 129
        43004 => X"78",  -- 120
        43005 => X"7A",  -- 122
        43006 => X"7D",  -- 125
        43007 => X"76",  -- 118
        43008 => X"69",  -- 105
        43009 => X"6E",  -- 110
        43010 => X"7C",  -- 124
        43011 => X"73",  -- 115
        43012 => X"79",  -- 121
        43013 => X"62",  -- 98
        43014 => X"35",  -- 53
        43015 => X"52",  -- 82
        43016 => X"9E",  -- 158
        43017 => X"BC",  -- 188
        43018 => X"CE",  -- 206
        43019 => X"D7",  -- 215
        43020 => X"CC",  -- 204
        43021 => X"C3",  -- 195
        43022 => X"CB",  -- 203
        43023 => X"C0",  -- 192
        43024 => X"82",  -- 130
        43025 => X"46",  -- 70
        43026 => X"75",  -- 117
        43027 => X"9A",  -- 154
        43028 => X"B6",  -- 182
        43029 => X"C6",  -- 198
        43030 => X"C7",  -- 199
        43031 => X"C6",  -- 198
        43032 => X"C6",  -- 198
        43033 => X"BF",  -- 191
        43034 => X"B4",  -- 180
        43035 => X"AB",  -- 171
        43036 => X"3E",  -- 62
        43037 => X"1E",  -- 30
        43038 => X"2B",  -- 43
        43039 => X"30",  -- 48
        43040 => X"6D",  -- 109
        43041 => X"92",  -- 146
        43042 => X"AC",  -- 172
        43043 => X"BA",  -- 186
        43044 => X"B3",  -- 179
        43045 => X"AF",  -- 175
        43046 => X"B3",  -- 179
        43047 => X"A4",  -- 164
        43048 => X"9B",  -- 155
        43049 => X"C0",  -- 192
        43050 => X"C2",  -- 194
        43051 => X"D2",  -- 210
        43052 => X"C0",  -- 192
        43053 => X"9A",  -- 154
        43054 => X"97",  -- 151
        43055 => X"80",  -- 128
        43056 => X"61",  -- 97
        43057 => X"63",  -- 99
        43058 => X"69",  -- 105
        43059 => X"64",  -- 100
        43060 => X"61",  -- 97
        43061 => X"67",  -- 103
        43062 => X"5F",  -- 95
        43063 => X"4F",  -- 79
        43064 => X"52",  -- 82
        43065 => X"4F",  -- 79
        43066 => X"4D",  -- 77
        43067 => X"4D",  -- 77
        43068 => X"51",  -- 81
        43069 => X"56",  -- 86
        43070 => X"5A",  -- 90
        43071 => X"5E",  -- 94
        43072 => X"5D",  -- 93
        43073 => X"58",  -- 88
        43074 => X"55",  -- 85
        43075 => X"56",  -- 86
        43076 => X"56",  -- 86
        43077 => X"52",  -- 82
        43078 => X"50",  -- 80
        43079 => X"51",  -- 81
        43080 => X"54",  -- 84
        43081 => X"51",  -- 81
        43082 => X"4F",  -- 79
        43083 => X"4F",  -- 79
        43084 => X"52",  -- 82
        43085 => X"55",  -- 85
        43086 => X"55",  -- 85
        43087 => X"53",  -- 83
        43088 => X"54",  -- 84
        43089 => X"52",  -- 82
        43090 => X"53",  -- 83
        43091 => X"55",  -- 85
        43092 => X"53",  -- 83
        43093 => X"4E",  -- 78
        43094 => X"4C",  -- 76
        43095 => X"4E",  -- 78
        43096 => X"45",  -- 69
        43097 => X"46",  -- 70
        43098 => X"47",  -- 71
        43099 => X"45",  -- 69
        43100 => X"43",  -- 67
        43101 => X"40",  -- 64
        43102 => X"3F",  -- 63
        43103 => X"40",  -- 64
        43104 => X"43",  -- 67
        43105 => X"43",  -- 67
        43106 => X"40",  -- 64
        43107 => X"3F",  -- 63
        43108 => X"44",  -- 68
        43109 => X"44",  -- 68
        43110 => X"50",  -- 80
        43111 => X"65",  -- 101
        43112 => X"77",  -- 119
        43113 => X"82",  -- 130
        43114 => X"92",  -- 146
        43115 => X"9D",  -- 157
        43116 => X"A9",  -- 169
        43117 => X"AF",  -- 175
        43118 => X"B0",  -- 176
        43119 => X"AE",  -- 174
        43120 => X"AA",  -- 170
        43121 => X"B1",  -- 177
        43122 => X"B6",  -- 182
        43123 => X"A3",  -- 163
        43124 => X"9E",  -- 158
        43125 => X"AD",  -- 173
        43126 => X"AF",  -- 175
        43127 => X"B5",  -- 181
        43128 => X"B4",  -- 180
        43129 => X"AF",  -- 175
        43130 => X"AE",  -- 174
        43131 => X"B0",  -- 176
        43132 => X"B1",  -- 177
        43133 => X"AF",  -- 175
        43134 => X"AE",  -- 174
        43135 => X"AD",  -- 173
        43136 => X"B1",  -- 177
        43137 => X"B6",  -- 182
        43138 => X"AE",  -- 174
        43139 => X"A4",  -- 164
        43140 => X"A7",  -- 167
        43141 => X"AA",  -- 170
        43142 => X"A7",  -- 167
        43143 => X"A3",  -- 163
        43144 => X"A2",  -- 162
        43145 => X"A1",  -- 161
        43146 => X"9F",  -- 159
        43147 => X"9E",  -- 158
        43148 => X"9E",  -- 158
        43149 => X"9E",  -- 158
        43150 => X"A2",  -- 162
        43151 => X"A6",  -- 166
        43152 => X"AF",  -- 175
        43153 => X"B3",  -- 179
        43154 => X"B0",  -- 176
        43155 => X"A9",  -- 169
        43156 => X"A8",  -- 168
        43157 => X"AF",  -- 175
        43158 => X"B2",  -- 178
        43159 => X"AE",  -- 174
        43160 => X"B1",  -- 177
        43161 => X"B3",  -- 179
        43162 => X"B0",  -- 176
        43163 => X"AB",  -- 171
        43164 => X"AC",  -- 172
        43165 => X"B7",  -- 183
        43166 => X"C1",  -- 193
        43167 => X"C6",  -- 198
        43168 => X"C5",  -- 197
        43169 => X"C8",  -- 200
        43170 => X"CB",  -- 203
        43171 => X"CD",  -- 205
        43172 => X"CD",  -- 205
        43173 => X"C8",  -- 200
        43174 => X"BC",  -- 188
        43175 => X"B0",  -- 176
        43176 => X"B1",  -- 177
        43177 => X"A8",  -- 168
        43178 => X"A5",  -- 165
        43179 => X"A5",  -- 165
        43180 => X"9E",  -- 158
        43181 => X"9C",  -- 156
        43182 => X"98",  -- 152
        43183 => X"8E",  -- 142
        43184 => X"89",  -- 137
        43185 => X"66",  -- 102
        43186 => X"6C",  -- 108
        43187 => X"55",  -- 85
        43188 => X"3B",  -- 59
        43189 => X"55",  -- 85
        43190 => X"67",  -- 103
        43191 => X"70",  -- 112
        43192 => X"68",  -- 104
        43193 => X"73",  -- 115
        43194 => X"81",  -- 129
        43195 => X"81",  -- 129
        43196 => X"74",  -- 116
        43197 => X"62",  -- 98
        43198 => X"58",  -- 88
        43199 => X"57",  -- 87
        43200 => X"61",  -- 97
        43201 => X"65",  -- 101
        43202 => X"6D",  -- 109
        43203 => X"73",  -- 115
        43204 => X"75",  -- 117
        43205 => X"73",  -- 115
        43206 => X"6B",  -- 107
        43207 => X"67",  -- 103
        43208 => X"66",  -- 102
        43209 => X"6E",  -- 110
        43210 => X"76",  -- 118
        43211 => X"78",  -- 120
        43212 => X"74",  -- 116
        43213 => X"6E",  -- 110
        43214 => X"6A",  -- 106
        43215 => X"6B",  -- 107
        43216 => X"62",  -- 98
        43217 => X"5D",  -- 93
        43218 => X"5B",  -- 91
        43219 => X"5A",  -- 90
        43220 => X"5A",  -- 90
        43221 => X"58",  -- 88
        43222 => X"53",  -- 83
        43223 => X"4F",  -- 79
        43224 => X"4E",  -- 78
        43225 => X"5A",  -- 90
        43226 => X"59",  -- 89
        43227 => X"58",  -- 88
        43228 => X"5B",  -- 91
        43229 => X"50",  -- 80
        43230 => X"51",  -- 81
        43231 => X"66",  -- 102
        43232 => X"8E",  -- 142
        43233 => X"75",  -- 117
        43234 => X"68",  -- 104
        43235 => X"54",  -- 84
        43236 => X"39",  -- 57
        43237 => X"22",  -- 34
        43238 => X"18",  -- 24
        43239 => X"2C",  -- 44
        43240 => X"5D",  -- 93
        43241 => X"69",  -- 105
        43242 => X"58",  -- 88
        43243 => X"51",  -- 81
        43244 => X"38",  -- 56
        43245 => X"16",  -- 22
        43246 => X"1C",  -- 28
        43247 => X"1D",  -- 29
        43248 => X"13",  -- 19
        43249 => X"44",  -- 68
        43250 => X"84",  -- 132
        43251 => X"91",  -- 145
        43252 => X"95",  -- 149
        43253 => X"8F",  -- 143
        43254 => X"6E",  -- 110
        43255 => X"6F",  -- 111
        43256 => X"53",  -- 83
        43257 => X"38",  -- 56
        43258 => X"22",  -- 34
        43259 => X"31",  -- 49
        43260 => X"47",  -- 71
        43261 => X"4B",  -- 75
        43262 => X"51",  -- 81
        43263 => X"66",  -- 102
        43264 => X"61",  -- 97
        43265 => X"5D",  -- 93
        43266 => X"59",  -- 89
        43267 => X"57",  -- 87
        43268 => X"60",  -- 96
        43269 => X"5E",  -- 94
        43270 => X"46",  -- 70
        43271 => X"3C",  -- 60
        43272 => X"24",  -- 36
        43273 => X"26",  -- 38
        43274 => X"24",  -- 36
        43275 => X"29",  -- 41
        43276 => X"36",  -- 54
        43277 => X"36",  -- 54
        43278 => X"2E",  -- 46
        43279 => X"2D",  -- 45
        43280 => X"32",  -- 50
        43281 => X"32",  -- 50
        43282 => X"36",  -- 54
        43283 => X"3B",  -- 59
        43284 => X"41",  -- 65
        43285 => X"47",  -- 71
        43286 => X"4F",  -- 79
        43287 => X"57",  -- 87
        43288 => X"5E",  -- 94
        43289 => X"60",  -- 96
        43290 => X"61",  -- 97
        43291 => X"5E",  -- 94
        43292 => X"5E",  -- 94
        43293 => X"60",  -- 96
        43294 => X"5E",  -- 94
        43295 => X"58",  -- 88
        43296 => X"61",  -- 97
        43297 => X"71",  -- 113
        43298 => X"72",  -- 114
        43299 => X"80",  -- 128
        43300 => X"82",  -- 130
        43301 => X"89",  -- 137
        43302 => X"7B",  -- 123
        43303 => X"7C",  -- 124
        43304 => X"69",  -- 105
        43305 => X"66",  -- 102
        43306 => X"60",  -- 96
        43307 => X"58",  -- 88
        43308 => X"53",  -- 83
        43309 => X"52",  -- 82
        43310 => X"51",  -- 81
        43311 => X"4F",  -- 79
        43312 => X"49",  -- 73
        43313 => X"40",  -- 64
        43314 => X"3A",  -- 58
        43315 => X"3A",  -- 58
        43316 => X"3C",  -- 60
        43317 => X"4E",  -- 78
        43318 => X"67",  -- 103
        43319 => X"70",  -- 112
        43320 => X"8B",  -- 139
        43321 => X"8A",  -- 138
        43322 => X"8C",  -- 140
        43323 => X"85",  -- 133
        43324 => X"7C",  -- 124
        43325 => X"80",  -- 128
        43326 => X"86",  -- 134
        43327 => X"81",  -- 129
        43328 => X"73",  -- 115
        43329 => X"70",  -- 112
        43330 => X"74",  -- 116
        43331 => X"6D",  -- 109
        43332 => X"8F",  -- 143
        43333 => X"9B",  -- 155
        43334 => X"7E",  -- 126
        43335 => X"9C",  -- 156
        43336 => X"BA",  -- 186
        43337 => X"C7",  -- 199
        43338 => X"C4",  -- 196
        43339 => X"BF",  -- 191
        43340 => X"B1",  -- 177
        43341 => X"B0",  -- 176
        43342 => X"B8",  -- 184
        43343 => X"96",  -- 150
        43344 => X"6F",  -- 111
        43345 => X"3E",  -- 62
        43346 => X"71",  -- 113
        43347 => X"81",  -- 129
        43348 => X"99",  -- 153
        43349 => X"B4",  -- 180
        43350 => X"BB",  -- 187
        43351 => X"BE",  -- 190
        43352 => X"AA",  -- 170
        43353 => X"AF",  -- 175
        43354 => X"A8",  -- 168
        43355 => X"AE",  -- 174
        43356 => X"3C",  -- 60
        43357 => X"19",  -- 25
        43358 => X"33",  -- 51
        43359 => X"30",  -- 48
        43360 => X"6F",  -- 111
        43361 => X"8C",  -- 140
        43362 => X"96",  -- 150
        43363 => X"B0",  -- 176
        43364 => X"C6",  -- 198
        43365 => X"B8",  -- 184
        43366 => X"AE",  -- 174
        43367 => X"B1",  -- 177
        43368 => X"A2",  -- 162
        43369 => X"B6",  -- 182
        43370 => X"C3",  -- 195
        43371 => X"CE",  -- 206
        43372 => X"C0",  -- 192
        43373 => X"96",  -- 150
        43374 => X"7C",  -- 124
        43375 => X"73",  -- 115
        43376 => X"5A",  -- 90
        43377 => X"59",  -- 89
        43378 => X"54",  -- 84
        43379 => X"64",  -- 100
        43380 => X"5F",  -- 95
        43381 => X"58",  -- 88
        43382 => X"64",  -- 100
        43383 => X"4D",  -- 77
        43384 => X"4A",  -- 74
        43385 => X"4C",  -- 76
        43386 => X"4F",  -- 79
        43387 => X"51",  -- 81
        43388 => X"52",  -- 82
        43389 => X"55",  -- 85
        43390 => X"57",  -- 87
        43391 => X"5A",  -- 90
        43392 => X"63",  -- 99
        43393 => X"59",  -- 89
        43394 => X"51",  -- 81
        43395 => X"52",  -- 82
        43396 => X"54",  -- 84
        43397 => X"52",  -- 82
        43398 => X"52",  -- 82
        43399 => X"54",  -- 84
        43400 => X"52",  -- 82
        43401 => X"51",  -- 81
        43402 => X"4F",  -- 79
        43403 => X"4E",  -- 78
        43404 => X"4F",  -- 79
        43405 => X"51",  -- 81
        43406 => X"50",  -- 80
        43407 => X"4E",  -- 78
        43408 => X"51",  -- 81
        43409 => X"4F",  -- 79
        43410 => X"51",  -- 81
        43411 => X"55",  -- 85
        43412 => X"53",  -- 83
        43413 => X"4D",  -- 77
        43414 => X"4B",  -- 75
        43415 => X"4D",  -- 77
        43416 => X"42",  -- 66
        43417 => X"44",  -- 68
        43418 => X"46",  -- 70
        43419 => X"46",  -- 70
        43420 => X"43",  -- 67
        43421 => X"3F",  -- 63
        43422 => X"3C",  -- 60
        43423 => X"3C",  -- 60
        43424 => X"45",  -- 69
        43425 => X"44",  -- 68
        43426 => X"40",  -- 64
        43427 => X"41",  -- 65
        43428 => X"46",  -- 70
        43429 => X"45",  -- 69
        43430 => X"51",  -- 81
        43431 => X"6A",  -- 106
        43432 => X"7A",  -- 122
        43433 => X"87",  -- 135
        43434 => X"95",  -- 149
        43435 => X"A0",  -- 160
        43436 => X"A6",  -- 166
        43437 => X"AA",  -- 170
        43438 => X"A9",  -- 169
        43439 => X"A6",  -- 166
        43440 => X"A6",  -- 166
        43441 => X"AA",  -- 170
        43442 => X"AE",  -- 174
        43443 => X"9E",  -- 158
        43444 => X"9A",  -- 154
        43445 => X"AC",  -- 172
        43446 => X"B0",  -- 176
        43447 => X"B5",  -- 181
        43448 => X"B9",  -- 185
        43449 => X"B3",  -- 179
        43450 => X"AB",  -- 171
        43451 => X"AA",  -- 170
        43452 => X"AC",  -- 172
        43453 => X"A4",  -- 164
        43454 => X"9D",  -- 157
        43455 => X"A2",  -- 162
        43456 => X"AF",  -- 175
        43457 => X"BB",  -- 187
        43458 => X"AE",  -- 174
        43459 => X"9D",  -- 157
        43460 => X"A5",  -- 165
        43461 => X"AA",  -- 170
        43462 => X"9E",  -- 158
        43463 => X"99",  -- 153
        43464 => X"98",  -- 152
        43465 => X"9B",  -- 155
        43466 => X"9E",  -- 158
        43467 => X"9A",  -- 154
        43468 => X"95",  -- 149
        43469 => X"97",  -- 151
        43470 => X"A2",  -- 162
        43471 => X"AB",  -- 171
        43472 => X"A8",  -- 168
        43473 => X"B2",  -- 178
        43474 => X"B5",  -- 181
        43475 => X"B0",  -- 176
        43476 => X"AC",  -- 172
        43477 => X"B1",  -- 177
        43478 => X"B6",  -- 182
        43479 => X"B5",  -- 181
        43480 => X"AB",  -- 171
        43481 => X"B4",  -- 180
        43482 => X"B7",  -- 183
        43483 => X"AF",  -- 175
        43484 => X"AA",  -- 170
        43485 => X"B1",  -- 177
        43486 => X"BE",  -- 190
        43487 => X"C7",  -- 199
        43488 => X"C3",  -- 195
        43489 => X"C5",  -- 197
        43490 => X"C8",  -- 200
        43491 => X"CC",  -- 204
        43492 => X"D1",  -- 209
        43493 => X"D0",  -- 208
        43494 => X"C6",  -- 198
        43495 => X"BA",  -- 186
        43496 => X"B7",  -- 183
        43497 => X"AB",  -- 171
        43498 => X"A6",  -- 166
        43499 => X"A5",  -- 165
        43500 => X"9F",  -- 159
        43501 => X"9C",  -- 156
        43502 => X"96",  -- 150
        43503 => X"8A",  -- 138
        43504 => X"72",  -- 114
        43505 => X"68",  -- 104
        43506 => X"45",  -- 69
        43507 => X"53",  -- 83
        43508 => X"55",  -- 85
        43509 => X"39",  -- 57
        43510 => X"53",  -- 83
        43511 => X"79",  -- 121
        43512 => X"84",  -- 132
        43513 => X"7A",  -- 122
        43514 => X"77",  -- 119
        43515 => X"76",  -- 118
        43516 => X"6A",  -- 106
        43517 => X"56",  -- 86
        43518 => X"50",  -- 80
        43519 => X"58",  -- 88
        43520 => X"66",  -- 102
        43521 => X"64",  -- 100
        43522 => X"67",  -- 103
        43523 => X"6C",  -- 108
        43524 => X"73",  -- 115
        43525 => X"75",  -- 117
        43526 => X"70",  -- 112
        43527 => X"6A",  -- 106
        43528 => X"6B",  -- 107
        43529 => X"71",  -- 113
        43530 => X"74",  -- 116
        43531 => X"74",  -- 116
        43532 => X"70",  -- 112
        43533 => X"6E",  -- 110
        43534 => X"70",  -- 112
        43535 => X"75",  -- 117
        43536 => X"6B",  -- 107
        43537 => X"62",  -- 98
        43538 => X"58",  -- 88
        43539 => X"53",  -- 83
        43540 => X"54",  -- 84
        43541 => X"54",  -- 84
        43542 => X"52",  -- 82
        43543 => X"4F",  -- 79
        43544 => X"56",  -- 86
        43545 => X"54",  -- 84
        43546 => X"53",  -- 83
        43547 => X"56",  -- 86
        43548 => X"57",  -- 87
        43549 => X"4F",  -- 79
        43550 => X"57",  -- 87
        43551 => X"6E",  -- 110
        43552 => X"8C",  -- 140
        43553 => X"79",  -- 121
        43554 => X"71",  -- 113
        43555 => X"53",  -- 83
        43556 => X"3D",  -- 61
        43557 => X"32",  -- 50
        43558 => X"18",  -- 24
        43559 => X"1A",  -- 26
        43560 => X"3B",  -- 59
        43561 => X"58",  -- 88
        43562 => X"4D",  -- 77
        43563 => X"20",  -- 32
        43564 => X"16",  -- 22
        43565 => X"14",  -- 20
        43566 => X"08",  -- 8
        43567 => X"21",  -- 33
        43568 => X"11",  -- 17
        43569 => X"20",  -- 32
        43570 => X"4A",  -- 74
        43571 => X"79",  -- 121
        43572 => X"8C",  -- 140
        43573 => X"8A",  -- 138
        43574 => X"83",  -- 131
        43575 => X"7A",  -- 122
        43576 => X"6F",  -- 111
        43577 => X"6B",  -- 107
        43578 => X"59",  -- 89
        43579 => X"55",  -- 85
        43580 => X"54",  -- 84
        43581 => X"57",  -- 87
        43582 => X"5E",  -- 94
        43583 => X"5A",  -- 90
        43584 => X"55",  -- 85
        43585 => X"62",  -- 98
        43586 => X"56",  -- 86
        43587 => X"63",  -- 99
        43588 => X"65",  -- 101
        43589 => X"4C",  -- 76
        43590 => X"42",  -- 66
        43591 => X"31",  -- 49
        43592 => X"2B",  -- 43
        43593 => X"2A",  -- 42
        43594 => X"2B",  -- 43
        43595 => X"2C",  -- 44
        43596 => X"2F",  -- 47
        43597 => X"31",  -- 49
        43598 => X"33",  -- 51
        43599 => X"32",  -- 50
        43600 => X"3B",  -- 59
        43601 => X"40",  -- 64
        43602 => X"48",  -- 72
        43603 => X"4D",  -- 77
        43604 => X"4D",  -- 77
        43605 => X"4D",  -- 77
        43606 => X"53",  -- 83
        43607 => X"5D",  -- 93
        43608 => X"5F",  -- 95
        43609 => X"61",  -- 97
        43610 => X"6A",  -- 106
        43611 => X"59",  -- 89
        43612 => X"5C",  -- 92
        43613 => X"55",  -- 85
        43614 => X"61",  -- 97
        43615 => X"5E",  -- 94
        43616 => X"74",  -- 116
        43617 => X"82",  -- 130
        43618 => X"79",  -- 121
        43619 => X"81",  -- 129
        43620 => X"85",  -- 133
        43621 => X"6A",  -- 106
        43622 => X"8A",  -- 138
        43623 => X"72",  -- 114
        43624 => X"6D",  -- 109
        43625 => X"79",  -- 121
        43626 => X"6A",  -- 106
        43627 => X"5D",  -- 93
        43628 => X"56",  -- 86
        43629 => X"50",  -- 80
        43630 => X"55",  -- 85
        43631 => X"52",  -- 82
        43632 => X"54",  -- 84
        43633 => X"38",  -- 56
        43634 => X"3B",  -- 59
        43635 => X"3B",  -- 59
        43636 => X"3F",  -- 63
        43637 => X"43",  -- 67
        43638 => X"65",  -- 101
        43639 => X"76",  -- 118
        43640 => X"85",  -- 133
        43641 => X"8C",  -- 140
        43642 => X"93",  -- 147
        43643 => X"92",  -- 146
        43644 => X"8B",  -- 139
        43645 => X"87",  -- 135
        43646 => X"89",  -- 137
        43647 => X"8E",  -- 142
        43648 => X"8B",  -- 139
        43649 => X"8E",  -- 142
        43650 => X"8D",  -- 141
        43651 => X"8C",  -- 140
        43652 => X"9A",  -- 154
        43653 => X"A5",  -- 165
        43654 => X"B1",  -- 177
        43655 => X"C0",  -- 192
        43656 => X"CD",  -- 205
        43657 => X"C2",  -- 194
        43658 => X"C2",  -- 194
        43659 => X"C6",  -- 198
        43660 => X"91",  -- 145
        43661 => X"96",  -- 150
        43662 => X"8B",  -- 139
        43663 => X"50",  -- 80
        43664 => X"22",  -- 34
        43665 => X"33",  -- 51
        43666 => X"3F",  -- 63
        43667 => X"4F",  -- 79
        43668 => X"95",  -- 149
        43669 => X"AE",  -- 174
        43670 => X"B7",  -- 183
        43671 => X"BB",  -- 187
        43672 => X"A6",  -- 166
        43673 => X"86",  -- 134
        43674 => X"8F",  -- 143
        43675 => X"75",  -- 117
        43676 => X"64",  -- 100
        43677 => X"2B",  -- 43
        43678 => X"3B",  -- 59
        43679 => X"46",  -- 70
        43680 => X"63",  -- 99
        43681 => X"84",  -- 132
        43682 => X"95",  -- 149
        43683 => X"7E",  -- 126
        43684 => X"B0",  -- 176
        43685 => X"B1",  -- 177
        43686 => X"BA",  -- 186
        43687 => X"B3",  -- 179
        43688 => X"AA",  -- 170
        43689 => X"A8",  -- 168
        43690 => X"C4",  -- 196
        43691 => X"C2",  -- 194
        43692 => X"AF",  -- 175
        43693 => X"95",  -- 149
        43694 => X"6D",  -- 109
        43695 => X"69",  -- 105
        43696 => X"5D",  -- 93
        43697 => X"52",  -- 82
        43698 => X"4A",  -- 74
        43699 => X"4B",  -- 75
        43700 => X"53",  -- 83
        43701 => X"58",  -- 88
        43702 => X"54",  -- 84
        43703 => X"4F",  -- 79
        43704 => X"49",  -- 73
        43705 => X"4D",  -- 77
        43706 => X"51",  -- 81
        43707 => X"50",  -- 80
        43708 => X"4D",  -- 77
        43709 => X"4E",  -- 78
        43710 => X"54",  -- 84
        43711 => X"5A",  -- 90
        43712 => X"5F",  -- 95
        43713 => X"5E",  -- 94
        43714 => X"55",  -- 85
        43715 => X"51",  -- 81
        43716 => X"56",  -- 86
        43717 => X"54",  -- 84
        43718 => X"4D",  -- 77
        43719 => X"4D",  -- 77
        43720 => X"52",  -- 82
        43721 => X"52",  -- 82
        43722 => X"50",  -- 80
        43723 => X"4E",  -- 78
        43724 => X"4C",  -- 76
        43725 => X"4B",  -- 75
        43726 => X"4C",  -- 76
        43727 => X"4D",  -- 77
        43728 => X"4E",  -- 78
        43729 => X"4E",  -- 78
        43730 => X"4C",  -- 76
        43731 => X"4B",  -- 75
        43732 => X"50",  -- 80
        43733 => X"54",  -- 84
        43734 => X"50",  -- 80
        43735 => X"48",  -- 72
        43736 => X"41",  -- 65
        43737 => X"44",  -- 68
        43738 => X"44",  -- 68
        43739 => X"43",  -- 67
        43740 => X"43",  -- 67
        43741 => X"44",  -- 68
        43742 => X"41",  -- 65
        43743 => X"3D",  -- 61
        43744 => X"41",  -- 65
        43745 => X"40",  -- 64
        43746 => X"42",  -- 66
        43747 => X"44",  -- 68
        43748 => X"41",  -- 65
        43749 => X"44",  -- 68
        43750 => X"57",  -- 87
        43751 => X"6F",  -- 111
        43752 => X"7D",  -- 125
        43753 => X"8E",  -- 142
        43754 => X"97",  -- 151
        43755 => X"9D",  -- 157
        43756 => X"A2",  -- 162
        43757 => X"A3",  -- 163
        43758 => X"A5",  -- 165
        43759 => X"AC",  -- 172
        43760 => X"9D",  -- 157
        43761 => X"B0",  -- 176
        43762 => X"B6",  -- 182
        43763 => X"A9",  -- 169
        43764 => X"A6",  -- 166
        43765 => X"B3",  -- 179
        43766 => X"B8",  -- 184
        43767 => X"B1",  -- 177
        43768 => X"AC",  -- 172
        43769 => X"B8",  -- 184
        43770 => X"AF",  -- 175
        43771 => X"AF",  -- 175
        43772 => X"A2",  -- 162
        43773 => X"AD",  -- 173
        43774 => X"A3",  -- 163
        43775 => X"A3",  -- 163
        43776 => X"A2",  -- 162
        43777 => X"BE",  -- 190
        43778 => X"A5",  -- 165
        43779 => X"9F",  -- 159
        43780 => X"A0",  -- 160
        43781 => X"A3",  -- 163
        43782 => X"96",  -- 150
        43783 => X"98",  -- 152
        43784 => X"98",  -- 152
        43785 => X"A3",  -- 163
        43786 => X"A8",  -- 168
        43787 => X"A0",  -- 160
        43788 => X"9A",  -- 154
        43789 => X"A1",  -- 161
        43790 => X"A4",  -- 164
        43791 => X"A2",  -- 162
        43792 => X"AE",  -- 174
        43793 => X"B1",  -- 177
        43794 => X"B5",  -- 181
        43795 => X"B6",  -- 182
        43796 => X"AF",  -- 175
        43797 => X"AD",  -- 173
        43798 => X"B6",  -- 182
        43799 => X"C2",  -- 194
        43800 => X"B8",  -- 184
        43801 => X"B1",  -- 177
        43802 => X"AB",  -- 171
        43803 => X"AD",  -- 173
        43804 => X"B1",  -- 177
        43805 => X"B4",  -- 180
        43806 => X"BA",  -- 186
        43807 => X"C1",  -- 193
        43808 => X"CA",  -- 202
        43809 => X"C7",  -- 199
        43810 => X"C7",  -- 199
        43811 => X"CC",  -- 204
        43812 => X"CF",  -- 207
        43813 => X"CC",  -- 204
        43814 => X"C8",  -- 200
        43815 => X"C5",  -- 197
        43816 => X"B9",  -- 185
        43817 => X"BA",  -- 186
        43818 => X"B6",  -- 182
        43819 => X"AC",  -- 172
        43820 => X"A1",  -- 161
        43821 => X"99",  -- 153
        43822 => X"8E",  -- 142
        43823 => X"85",  -- 133
        43824 => X"88",  -- 136
        43825 => X"71",  -- 113
        43826 => X"4D",  -- 77
        43827 => X"3D",  -- 61
        43828 => X"3E",  -- 62
        43829 => X"3C",  -- 60
        43830 => X"4C",  -- 76
        43831 => X"71",  -- 113
        43832 => X"7D",  -- 125
        43833 => X"85",  -- 133
        43834 => X"81",  -- 129
        43835 => X"7D",  -- 125
        43836 => X"77",  -- 119
        43837 => X"4D",  -- 77
        43838 => X"30",  -- 48
        43839 => X"3F",  -- 63
        43840 => X"6E",  -- 110
        43841 => X"68",  -- 104
        43842 => X"64",  -- 100
        43843 => X"64",  -- 100
        43844 => X"69",  -- 105
        43845 => X"70",  -- 112
        43846 => X"71",  -- 113
        43847 => X"70",  -- 112
        43848 => X"77",  -- 119
        43849 => X"7A",  -- 122
        43850 => X"7B",  -- 123
        43851 => X"78",  -- 120
        43852 => X"73",  -- 115
        43853 => X"70",  -- 112
        43854 => X"6F",  -- 111
        43855 => X"72",  -- 114
        43856 => X"72",  -- 114
        43857 => X"69",  -- 105
        43858 => X"5D",  -- 93
        43859 => X"57",  -- 87
        43860 => X"55",  -- 85
        43861 => X"53",  -- 83
        43862 => X"51",  -- 81
        43863 => X"50",  -- 80
        43864 => X"51",  -- 81
        43865 => X"53",  -- 83
        43866 => X"55",  -- 85
        43867 => X"56",  -- 86
        43868 => X"55",  -- 85
        43869 => X"4F",  -- 79
        43870 => X"5D",  -- 93
        43871 => X"79",  -- 121
        43872 => X"88",  -- 136
        43873 => X"74",  -- 116
        43874 => X"71",  -- 113
        43875 => X"57",  -- 87
        43876 => X"4B",  -- 75
        43877 => X"2A",  -- 42
        43878 => X"1D",  -- 29
        43879 => X"1C",  -- 28
        43880 => X"32",  -- 50
        43881 => X"53",  -- 83
        43882 => X"53",  -- 83
        43883 => X"22",  -- 34
        43884 => X"0D",  -- 13
        43885 => X"0E",  -- 14
        43886 => X"03",  -- 3
        43887 => X"0E",  -- 14
        43888 => X"16",  -- 22
        43889 => X"15",  -- 21
        43890 => X"2B",  -- 43
        43891 => X"59",  -- 89
        43892 => X"81",  -- 129
        43893 => X"8A",  -- 138
        43894 => X"82",  -- 130
        43895 => X"7E",  -- 126
        43896 => X"79",  -- 121
        43897 => X"6A",  -- 106
        43898 => X"63",  -- 99
        43899 => X"61",  -- 97
        43900 => X"5D",  -- 93
        43901 => X"59",  -- 89
        43902 => X"5A",  -- 90
        43903 => X"62",  -- 98
        43904 => X"63",  -- 99
        43905 => X"68",  -- 104
        43906 => X"61",  -- 97
        43907 => X"64",  -- 100
        43908 => X"66",  -- 102
        43909 => X"52",  -- 82
        43910 => X"43",  -- 67
        43911 => X"39",  -- 57
        43912 => X"2A",  -- 42
        43913 => X"2B",  -- 43
        43914 => X"2D",  -- 45
        43915 => X"30",  -- 48
        43916 => X"31",  -- 49
        43917 => X"30",  -- 48
        43918 => X"38",  -- 56
        43919 => X"40",  -- 64
        43920 => X"4D",  -- 77
        43921 => X"44",  -- 68
        43922 => X"42",  -- 66
        43923 => X"49",  -- 73
        43924 => X"56",  -- 86
        43925 => X"5D",  -- 93
        43926 => X"5D",  -- 93
        43927 => X"5E",  -- 94
        43928 => X"66",  -- 102
        43929 => X"69",  -- 105
        43930 => X"6C",  -- 108
        43931 => X"6E",  -- 110
        43932 => X"67",  -- 103
        43933 => X"6D",  -- 109
        43934 => X"70",  -- 112
        43935 => X"6C",  -- 108
        43936 => X"70",  -- 112
        43937 => X"73",  -- 115
        43938 => X"83",  -- 131
        43939 => X"85",  -- 133
        43940 => X"87",  -- 135
        43941 => X"6E",  -- 110
        43942 => X"76",  -- 118
        43943 => X"7D",  -- 125
        43944 => X"7E",  -- 126
        43945 => X"85",  -- 133
        43946 => X"6D",  -- 109
        43947 => X"60",  -- 96
        43948 => X"60",  -- 96
        43949 => X"5C",  -- 92
        43950 => X"57",  -- 87
        43951 => X"47",  -- 71
        43952 => X"4B",  -- 75
        43953 => X"4F",  -- 79
        43954 => X"46",  -- 70
        43955 => X"3B",  -- 59
        43956 => X"58",  -- 88
        43957 => X"4C",  -- 76
        43958 => X"51",  -- 81
        43959 => X"6E",  -- 110
        43960 => X"87",  -- 135
        43961 => X"87",  -- 135
        43962 => X"88",  -- 136
        43963 => X"88",  -- 136
        43964 => X"89",  -- 137
        43965 => X"8F",  -- 143
        43966 => X"97",  -- 151
        43967 => X"9D",  -- 157
        43968 => X"92",  -- 146
        43969 => X"84",  -- 132
        43970 => X"7F",  -- 127
        43971 => X"87",  -- 135
        43972 => X"8A",  -- 138
        43973 => X"9D",  -- 157
        43974 => X"B8",  -- 184
        43975 => X"B3",  -- 179
        43976 => X"C3",  -- 195
        43977 => X"BD",  -- 189
        43978 => X"C5",  -- 197
        43979 => X"B1",  -- 177
        43980 => X"7B",  -- 123
        43981 => X"71",  -- 113
        43982 => X"5C",  -- 92
        43983 => X"2C",  -- 44
        43984 => X"30",  -- 48
        43985 => X"31",  -- 49
        43986 => X"35",  -- 53
        43987 => X"4E",  -- 78
        43988 => X"94",  -- 148
        43989 => X"AC",  -- 172
        43990 => X"B6",  -- 182
        43991 => X"C1",  -- 193
        43992 => X"A0",  -- 160
        43993 => X"76",  -- 118
        43994 => X"65",  -- 101
        43995 => X"5D",  -- 93
        43996 => X"53",  -- 83
        43997 => X"37",  -- 55
        43998 => X"41",  -- 65
        43999 => X"52",  -- 82
        44000 => X"6D",  -- 109
        44001 => X"7C",  -- 124
        44002 => X"89",  -- 137
        44003 => X"8F",  -- 143
        44004 => X"9F",  -- 159
        44005 => X"AE",  -- 174
        44006 => X"B8",  -- 184
        44007 => X"BA",  -- 186
        44008 => X"B6",  -- 182
        44009 => X"A9",  -- 169
        44010 => X"BF",  -- 191
        44011 => X"CA",  -- 202
        44012 => X"AE",  -- 174
        44013 => X"8B",  -- 139
        44014 => X"6A",  -- 106
        44015 => X"56",  -- 86
        44016 => X"56",  -- 86
        44017 => X"50",  -- 80
        44018 => X"48",  -- 72
        44019 => X"4A",  -- 74
        44020 => X"4F",  -- 79
        44021 => X"54",  -- 84
        44022 => X"51",  -- 81
        44023 => X"4C",  -- 76
        44024 => X"46",  -- 70
        44025 => X"4B",  -- 75
        44026 => X"4F",  -- 79
        44027 => X"4F",  -- 79
        44028 => X"4D",  -- 77
        44029 => X"4E",  -- 78
        44030 => X"53",  -- 83
        44031 => X"57",  -- 87
        44032 => X"5A",  -- 90
        44033 => X"5B",  -- 91
        44034 => X"53",  -- 83
        44035 => X"4F",  -- 79
        44036 => X"53",  -- 83
        44037 => X"51",  -- 81
        44038 => X"4B",  -- 75
        44039 => X"4D",  -- 77
        44040 => X"51",  -- 81
        44041 => X"51",  -- 81
        44042 => X"50",  -- 80
        44043 => X"4D",  -- 77
        44044 => X"4A",  -- 74
        44045 => X"49",  -- 73
        44046 => X"49",  -- 73
        44047 => X"4A",  -- 74
        44048 => X"4C",  -- 76
        44049 => X"4C",  -- 76
        44050 => X"4A",  -- 74
        44051 => X"4A",  -- 74
        44052 => X"4E",  -- 78
        44053 => X"52",  -- 82
        44054 => X"4E",  -- 78
        44055 => X"47",  -- 71
        44056 => X"42",  -- 66
        44057 => X"44",  -- 68
        44058 => X"43",  -- 67
        44059 => X"41",  -- 65
        44060 => X"42",  -- 66
        44061 => X"44",  -- 68
        44062 => X"43",  -- 67
        44063 => X"3F",  -- 63
        44064 => X"42",  -- 66
        44065 => X"41",  -- 65
        44066 => X"43",  -- 67
        44067 => X"45",  -- 69
        44068 => X"41",  -- 65
        44069 => X"44",  -- 68
        44070 => X"56",  -- 86
        44071 => X"6D",  -- 109
        44072 => X"7F",  -- 127
        44073 => X"90",  -- 144
        44074 => X"9C",  -- 156
        44075 => X"9F",  -- 159
        44076 => X"A4",  -- 164
        44077 => X"A4",  -- 164
        44078 => X"9E",  -- 158
        44079 => X"A0",  -- 160
        44080 => X"9E",  -- 158
        44081 => X"A6",  -- 166
        44082 => X"AA",  -- 170
        44083 => X"A9",  -- 169
        44084 => X"AA",  -- 170
        44085 => X"AF",  -- 175
        44086 => X"AD",  -- 173
        44087 => X"A7",  -- 167
        44088 => X"B0",  -- 176
        44089 => X"B4",  -- 180
        44090 => X"AE",  -- 174
        44091 => X"AA",  -- 170
        44092 => X"A6",  -- 166
        44093 => X"AF",  -- 175
        44094 => X"A7",  -- 167
        44095 => X"A0",  -- 160
        44096 => X"9C",  -- 156
        44097 => X"B2",  -- 178
        44098 => X"9B",  -- 155
        44099 => X"9D",  -- 157
        44100 => X"A0",  -- 160
        44101 => X"9E",  -- 158
        44102 => X"90",  -- 144
        44103 => X"93",  -- 147
        44104 => X"96",  -- 150
        44105 => X"9C",  -- 156
        44106 => X"9D",  -- 157
        44107 => X"96",  -- 150
        44108 => X"96",  -- 150
        44109 => X"A2",  -- 162
        44110 => X"AA",  -- 170
        44111 => X"AB",  -- 171
        44112 => X"AB",  -- 171
        44113 => X"AD",  -- 173
        44114 => X"B3",  -- 179
        44115 => X"B6",  -- 182
        44116 => X"B2",  -- 178
        44117 => X"AD",  -- 173
        44118 => X"AE",  -- 174
        44119 => X"B3",  -- 179
        44120 => X"B6",  -- 182
        44121 => X"B0",  -- 176
        44122 => X"AB",  -- 171
        44123 => X"AF",  -- 175
        44124 => X"B4",  -- 180
        44125 => X"B9",  -- 185
        44126 => X"BD",  -- 189
        44127 => X"C0",  -- 192
        44128 => X"CB",  -- 203
        44129 => X"C8",  -- 200
        44130 => X"C6",  -- 198
        44131 => X"C8",  -- 200
        44132 => X"CC",  -- 204
        44133 => X"CE",  -- 206
        44134 => X"CA",  -- 202
        44135 => X"C5",  -- 197
        44136 => X"BD",  -- 189
        44137 => X"BC",  -- 188
        44138 => X"B7",  -- 183
        44139 => X"B0",  -- 176
        44140 => X"A9",  -- 169
        44141 => X"9F",  -- 159
        44142 => X"8E",  -- 142
        44143 => X"7F",  -- 127
        44144 => X"61",  -- 97
        44145 => X"6D",  -- 109
        44146 => X"5F",  -- 95
        44147 => X"3F",  -- 63
        44148 => X"32",  -- 50
        44149 => X"3C",  -- 60
        44150 => X"49",  -- 73
        44151 => X"4F",  -- 79
        44152 => X"7A",  -- 122
        44153 => X"8C",  -- 140
        44154 => X"8D",  -- 141
        44155 => X"85",  -- 133
        44156 => X"82",  -- 130
        44157 => X"60",  -- 96
        44158 => X"3A",  -- 58
        44159 => X"35",  -- 53
        44160 => X"71",  -- 113
        44161 => X"6A",  -- 106
        44162 => X"64",  -- 100
        44163 => X"64",  -- 100
        44164 => X"67",  -- 103
        44165 => X"6F",  -- 111
        44166 => X"75",  -- 117
        44167 => X"77",  -- 119
        44168 => X"7C",  -- 124
        44169 => X"7C",  -- 124
        44170 => X"7C",  -- 124
        44171 => X"78",  -- 120
        44172 => X"73",  -- 115
        44173 => X"70",  -- 112
        44174 => X"70",  -- 112
        44175 => X"70",  -- 112
        44176 => X"72",  -- 114
        44177 => X"6B",  -- 107
        44178 => X"61",  -- 97
        44179 => X"59",  -- 89
        44180 => X"54",  -- 84
        44181 => X"53",  -- 83
        44182 => X"51",  -- 81
        44183 => X"51",  -- 81
        44184 => X"51",  -- 81
        44185 => X"59",  -- 89
        44186 => X"5B",  -- 91
        44187 => X"5B",  -- 91
        44188 => X"58",  -- 88
        44189 => X"51",  -- 81
        44190 => X"62",  -- 98
        44191 => X"80",  -- 128
        44192 => X"82",  -- 130
        44193 => X"71",  -- 113
        44194 => X"6F",  -- 111
        44195 => X"5E",  -- 94
        44196 => X"59",  -- 89
        44197 => X"25",  -- 37
        44198 => X"26",  -- 38
        44199 => X"21",  -- 33
        44200 => X"21",  -- 33
        44201 => X"42",  -- 66
        44202 => X"51",  -- 81
        44203 => X"24",  -- 36
        44204 => X"06",  -- 6
        44205 => X"0C",  -- 12
        44206 => X"0A",  -- 10
        44207 => X"09",  -- 9
        44208 => X"14",  -- 20
        44209 => X"0E",  -- 14
        44210 => X"0F",  -- 15
        44211 => X"32",  -- 50
        44212 => X"60",  -- 96
        44213 => X"6E",  -- 110
        44214 => X"74",  -- 116
        44215 => X"86",  -- 134
        44216 => X"86",  -- 134
        44217 => X"69",  -- 105
        44218 => X"66",  -- 102
        44219 => X"59",  -- 89
        44220 => X"51",  -- 81
        44221 => X"5B",  -- 91
        44222 => X"5D",  -- 93
        44223 => X"6B",  -- 107
        44224 => X"65",  -- 101
        44225 => X"65",  -- 101
        44226 => X"67",  -- 103
        44227 => X"63",  -- 99
        44228 => X"5F",  -- 95
        44229 => X"4F",  -- 79
        44230 => X"37",  -- 55
        44231 => X"37",  -- 55
        44232 => X"31",  -- 49
        44233 => X"2E",  -- 46
        44234 => X"31",  -- 49
        44235 => X"36",  -- 54
        44236 => X"30",  -- 48
        44237 => X"2B",  -- 43
        44238 => X"36",  -- 54
        44239 => X"48",  -- 72
        44240 => X"50",  -- 80
        44241 => X"4E",  -- 78
        44242 => X"4F",  -- 79
        44243 => X"55",  -- 85
        44244 => X"5C",  -- 92
        44245 => X"62",  -- 98
        44246 => X"69",  -- 105
        44247 => X"71",  -- 113
        44248 => X"6F",  -- 111
        44249 => X"6D",  -- 109
        44250 => X"6D",  -- 109
        44251 => X"7D",  -- 125
        44252 => X"6B",  -- 107
        44253 => X"7B",  -- 123
        44254 => X"77",  -- 119
        44255 => X"6E",  -- 110
        44256 => X"7C",  -- 124
        44257 => X"6B",  -- 107
        44258 => X"83",  -- 131
        44259 => X"80",  -- 128
        44260 => X"95",  -- 149
        44261 => X"8C",  -- 140
        44262 => X"6D",  -- 109
        44263 => X"84",  -- 132
        44264 => X"75",  -- 117
        44265 => X"8C",  -- 140
        44266 => X"7D",  -- 125
        44267 => X"6B",  -- 107
        44268 => X"61",  -- 97
        44269 => X"5C",  -- 92
        44270 => X"5E",  -- 94
        44271 => X"53",  -- 83
        44272 => X"44",  -- 68
        44273 => X"54",  -- 84
        44274 => X"53",  -- 83
        44275 => X"4A",  -- 74
        44276 => X"62",  -- 98
        44277 => X"52",  -- 82
        44278 => X"4F",  -- 79
        44279 => X"63",  -- 99
        44280 => X"84",  -- 132
        44281 => X"83",  -- 131
        44282 => X"84",  -- 132
        44283 => X"85",  -- 133
        44284 => X"88",  -- 136
        44285 => X"8B",  -- 139
        44286 => X"8E",  -- 142
        44287 => X"8E",  -- 142
        44288 => X"92",  -- 146
        44289 => X"89",  -- 137
        44290 => X"76",  -- 118
        44291 => X"83",  -- 131
        44292 => X"8E",  -- 142
        44293 => X"9D",  -- 157
        44294 => X"BE",  -- 190
        44295 => X"C1",  -- 193
        44296 => X"C3",  -- 195
        44297 => X"B6",  -- 182
        44298 => X"BB",  -- 187
        44299 => X"83",  -- 131
        44300 => X"52",  -- 82
        44301 => X"47",  -- 71
        44302 => X"3B",  -- 59
        44303 => X"2D",  -- 45
        44304 => X"3A",  -- 58
        44305 => X"29",  -- 41
        44306 => X"26",  -- 38
        44307 => X"44",  -- 68
        44308 => X"8B",  -- 139
        44309 => X"A2",  -- 162
        44310 => X"B3",  -- 179
        44311 => X"C3",  -- 195
        44312 => X"AF",  -- 175
        44313 => X"79",  -- 121
        44314 => X"4C",  -- 76
        44315 => X"50",  -- 80
        44316 => X"4D",  -- 77
        44317 => X"4A",  -- 74
        44318 => X"4B",  -- 75
        44319 => X"5F",  -- 95
        44320 => X"78",  -- 120
        44321 => X"76",  -- 118
        44322 => X"7A",  -- 122
        44323 => X"9C",  -- 156
        44324 => X"90",  -- 144
        44325 => X"AC",  -- 172
        44326 => X"B4",  -- 180
        44327 => X"BF",  -- 191
        44328 => X"BC",  -- 188
        44329 => X"A9",  -- 169
        44330 => X"B0",  -- 176
        44331 => X"C9",  -- 201
        44332 => X"B6",  -- 182
        44333 => X"8A",  -- 138
        44334 => X"6B",  -- 107
        44335 => X"4C",  -- 76
        44336 => X"4F",  -- 79
        44337 => X"4A",  -- 74
        44338 => X"46",  -- 70
        44339 => X"46",  -- 70
        44340 => X"49",  -- 73
        44341 => X"4C",  -- 76
        44342 => X"4B",  -- 75
        44343 => X"48",  -- 72
        44344 => X"42",  -- 66
        44345 => X"46",  -- 70
        44346 => X"4C",  -- 76
        44347 => X"4E",  -- 78
        44348 => X"4F",  -- 79
        44349 => X"4F",  -- 79
        44350 => X"52",  -- 82
        44351 => X"54",  -- 84
        44352 => X"53",  -- 83
        44353 => X"56",  -- 86
        44354 => X"51",  -- 81
        44355 => X"4D",  -- 77
        44356 => X"50",  -- 80
        44357 => X"4D",  -- 77
        44358 => X"49",  -- 73
        44359 => X"4D",  -- 77
        44360 => X"50",  -- 80
        44361 => X"50",  -- 80
        44362 => X"4F",  -- 79
        44363 => X"4C",  -- 76
        44364 => X"48",  -- 72
        44365 => X"46",  -- 70
        44366 => X"45",  -- 69
        44367 => X"46",  -- 70
        44368 => X"49",  -- 73
        44369 => X"48",  -- 72
        44370 => X"47",  -- 71
        44371 => X"48",  -- 72
        44372 => X"4C",  -- 76
        44373 => X"4F",  -- 79
        44374 => X"4C",  -- 76
        44375 => X"46",  -- 70
        44376 => X"42",  -- 66
        44377 => X"43",  -- 67
        44378 => X"42",  -- 66
        44379 => X"3F",  -- 63
        44380 => X"41",  -- 65
        44381 => X"44",  -- 68
        44382 => X"44",  -- 68
        44383 => X"43",  -- 67
        44384 => X"43",  -- 67
        44385 => X"42",  -- 66
        44386 => X"44",  -- 68
        44387 => X"44",  -- 68
        44388 => X"41",  -- 65
        44389 => X"45",  -- 69
        44390 => X"56",  -- 86
        44391 => X"6B",  -- 107
        44392 => X"7F",  -- 127
        44393 => X"94",  -- 148
        44394 => X"A0",  -- 160
        44395 => X"A0",  -- 160
        44396 => X"A7",  -- 167
        44397 => X"A6",  -- 166
        44398 => X"9A",  -- 154
        44399 => X"92",  -- 146
        44400 => X"97",  -- 151
        44401 => X"93",  -- 147
        44402 => X"97",  -- 151
        44403 => X"A3",  -- 163
        44404 => X"AD",  -- 173
        44405 => X"A9",  -- 169
        44406 => X"A3",  -- 163
        44407 => X"9D",  -- 157
        44408 => X"AE",  -- 174
        44409 => X"AA",  -- 170
        44410 => X"A7",  -- 167
        44411 => X"9F",  -- 159
        44412 => X"A6",  -- 166
        44413 => X"A6",  -- 166
        44414 => X"A0",  -- 160
        44415 => X"93",  -- 147
        44416 => X"9A",  -- 154
        44417 => X"AE",  -- 174
        44418 => X"9C",  -- 156
        44419 => X"A3",  -- 163
        44420 => X"A6",  -- 166
        44421 => X"A3",  -- 163
        44422 => X"95",  -- 149
        44423 => X"94",  -- 148
        44424 => X"90",  -- 144
        44425 => X"93",  -- 147
        44426 => X"93",  -- 147
        44427 => X"91",  -- 145
        44428 => X"97",  -- 151
        44429 => X"A5",  -- 165
        44430 => X"AD",  -- 173
        44431 => X"B0",  -- 176
        44432 => X"AC",  -- 172
        44433 => X"AD",  -- 173
        44434 => X"B0",  -- 176
        44435 => X"B4",  -- 180
        44436 => X"B2",  -- 178
        44437 => X"AE",  -- 174
        44438 => X"AC",  -- 172
        44439 => X"AD",  -- 173
        44440 => X"B2",  -- 178
        44441 => X"AC",  -- 172
        44442 => X"AB",  -- 171
        44443 => X"B1",  -- 177
        44444 => X"B7",  -- 183
        44445 => X"BA",  -- 186
        44446 => X"BC",  -- 188
        44447 => X"BE",  -- 190
        44448 => X"CA",  -- 202
        44449 => X"CA",  -- 202
        44450 => X"C6",  -- 198
        44451 => X"C2",  -- 194
        44452 => X"C6",  -- 198
        44453 => X"CD",  -- 205
        44454 => X"CC",  -- 204
        44455 => X"C7",  -- 199
        44456 => X"C0",  -- 192
        44457 => X"BC",  -- 188
        44458 => X"B6",  -- 182
        44459 => X"B2",  -- 178
        44460 => X"AF",  -- 175
        44461 => X"A5",  -- 165
        44462 => X"90",  -- 144
        44463 => X"7F",  -- 127
        44464 => X"6C",  -- 108
        44465 => X"51",  -- 81
        44466 => X"43",  -- 67
        44467 => X"41",  -- 65
        44468 => X"36",  -- 54
        44469 => X"2F",  -- 47
        44470 => X"3C",  -- 60
        44471 => X"4E",  -- 78
        44472 => X"60",  -- 96
        44473 => X"88",  -- 136
        44474 => X"9A",  -- 154
        44475 => X"92",  -- 146
        44476 => X"8B",  -- 139
        44477 => X"71",  -- 113
        44478 => X"4D",  -- 77
        44479 => X"3F",  -- 63
        44480 => X"6B",  -- 107
        44481 => X"6A",  -- 106
        44482 => X"6A",  -- 106
        44483 => X"6E",  -- 110
        44484 => X"72",  -- 114
        44485 => X"77",  -- 119
        44486 => X"7A",  -- 122
        44487 => X"7C",  -- 124
        44488 => X"78",  -- 120
        44489 => X"77",  -- 119
        44490 => X"76",  -- 118
        44491 => X"74",  -- 116
        44492 => X"72",  -- 114
        44493 => X"70",  -- 112
        44494 => X"70",  -- 112
        44495 => X"6E",  -- 110
        44496 => X"6C",  -- 108
        44497 => X"68",  -- 104
        44498 => X"5F",  -- 95
        44499 => X"58",  -- 88
        44500 => X"53",  -- 83
        44501 => X"51",  -- 81
        44502 => X"52",  -- 82
        44503 => X"52",  -- 82
        44504 => X"57",  -- 87
        44505 => X"5F",  -- 95
        44506 => X"62",  -- 98
        44507 => X"61",  -- 97
        44508 => X"5D",  -- 93
        44509 => X"55",  -- 85
        44510 => X"61",  -- 97
        44511 => X"7C",  -- 124
        44512 => X"78",  -- 120
        44513 => X"77",  -- 119
        44514 => X"6B",  -- 107
        44515 => X"67",  -- 103
        44516 => X"5B",  -- 91
        44517 => X"30",  -- 48
        44518 => X"33",  -- 51
        44519 => X"29",  -- 41
        44520 => X"1F",  -- 31
        44521 => X"36",  -- 54
        44522 => X"4F",  -- 79
        44523 => X"31",  -- 49
        44524 => X"0C",  -- 12
        44525 => X"0C",  -- 12
        44526 => X"0E",  -- 14
        44527 => X"0B",  -- 11
        44528 => X"04",  -- 4
        44529 => X"09",  -- 9
        44530 => X"06",  -- 6
        44531 => X"13",  -- 19
        44532 => X"2C",  -- 44
        44533 => X"33",  -- 51
        44534 => X"4B",  -- 75
        44535 => X"7E",  -- 126
        44536 => X"78",  -- 120
        44537 => X"52",  -- 82
        44538 => X"52",  -- 82
        44539 => X"3F",  -- 63
        44540 => X"40",  -- 64
        44541 => X"5F",  -- 95
        44542 => X"5F",  -- 95
        44543 => X"6A",  -- 106
        44544 => X"5E",  -- 94
        44545 => X"5D",  -- 93
        44546 => X"6C",  -- 108
        44547 => X"60",  -- 96
        44548 => X"55",  -- 85
        44549 => X"45",  -- 69
        44550 => X"28",  -- 40
        44551 => X"34",  -- 52
        44552 => X"3E",  -- 62
        44553 => X"37",  -- 55
        44554 => X"36",  -- 54
        44555 => X"38",  -- 56
        44556 => X"30",  -- 48
        44557 => X"25",  -- 37
        44558 => X"2D",  -- 45
        44559 => X"40",  -- 64
        44560 => X"48",  -- 72
        44561 => X"4D",  -- 77
        44562 => X"54",  -- 84
        44563 => X"5C",  -- 92
        44564 => X"61",  -- 97
        44565 => X"65",  -- 101
        44566 => X"6E",  -- 110
        44567 => X"77",  -- 119
        44568 => X"74",  -- 116
        44569 => X"6F",  -- 111
        44570 => X"73",  -- 115
        44571 => X"7F",  -- 127
        44572 => X"6E",  -- 110
        44573 => X"78",  -- 120
        44574 => X"77",  -- 119
        44575 => X"6B",  -- 107
        44576 => X"77",  -- 119
        44577 => X"6B",  -- 107
        44578 => X"78",  -- 120
        44579 => X"76",  -- 118
        44580 => X"92",  -- 146
        44581 => X"96",  -- 150
        44582 => X"6F",  -- 111
        44583 => X"85",  -- 133
        44584 => X"72",  -- 114
        44585 => X"8E",  -- 142
        44586 => X"85",  -- 133
        44587 => X"6E",  -- 110
        44588 => X"5F",  -- 95
        44589 => X"5B",  -- 91
        44590 => X"62",  -- 98
        44591 => X"5B",  -- 91
        44592 => X"47",  -- 71
        44593 => X"48",  -- 72
        44594 => X"5C",  -- 92
        44595 => X"5A",  -- 90
        44596 => X"57",  -- 87
        44597 => X"51",  -- 81
        44598 => X"63",  -- 99
        44599 => X"61",  -- 97
        44600 => X"79",  -- 121
        44601 => X"81",  -- 129
        44602 => X"8A",  -- 138
        44603 => X"90",  -- 144
        44604 => X"8F",  -- 143
        44605 => X"89",  -- 137
        44606 => X"7E",  -- 126
        44607 => X"75",  -- 117
        44608 => X"80",  -- 128
        44609 => X"9B",  -- 155
        44610 => X"83",  -- 131
        44611 => X"7B",  -- 123
        44612 => X"71",  -- 113
        44613 => X"5B",  -- 91
        44614 => X"7C",  -- 124
        44615 => X"A8",  -- 168
        44616 => X"96",  -- 150
        44617 => X"85",  -- 133
        44618 => X"86",  -- 134
        44619 => X"40",  -- 64
        44620 => X"25",  -- 37
        44621 => X"24",  -- 36
        44622 => X"24",  -- 36
        44623 => X"2E",  -- 46
        44624 => X"32",  -- 50
        44625 => X"1D",  -- 29
        44626 => X"19",  -- 25
        44627 => X"32",  -- 50
        44628 => X"76",  -- 118
        44629 => X"94",  -- 148
        44630 => X"AD",  -- 173
        44631 => X"B8",  -- 184
        44632 => X"AF",  -- 175
        44633 => X"7C",  -- 124
        44634 => X"4D",  -- 77
        44635 => X"51",  -- 81
        44636 => X"59",  -- 89
        44637 => X"5A",  -- 90
        44638 => X"5A",  -- 90
        44639 => X"6D",  -- 109
        44640 => X"7E",  -- 126
        44641 => X"7D",  -- 125
        44642 => X"77",  -- 119
        44643 => X"96",  -- 150
        44644 => X"91",  -- 145
        44645 => X"AE",  -- 174
        44646 => X"AE",  -- 174
        44647 => X"BB",  -- 187
        44648 => X"C4",  -- 196
        44649 => X"B5",  -- 181
        44650 => X"A1",  -- 161
        44651 => X"BC",  -- 188
        44652 => X"BF",  -- 191
        44653 => X"8E",  -- 142
        44654 => X"68",  -- 104
        44655 => X"4C",  -- 76
        44656 => X"4A",  -- 74
        44657 => X"47",  -- 71
        44658 => X"45",  -- 69
        44659 => X"44",  -- 68
        44660 => X"45",  -- 69
        44661 => X"47",  -- 71
        44662 => X"47",  -- 71
        44663 => X"46",  -- 70
        44664 => X"40",  -- 64
        44665 => X"44",  -- 68
        44666 => X"4A",  -- 74
        44667 => X"4E",  -- 78
        44668 => X"50",  -- 80
        44669 => X"50",  -- 80
        44670 => X"50",  -- 80
        44671 => X"50",  -- 80
        44672 => X"4C",  -- 76
        44673 => X"51",  -- 81
        44674 => X"4E",  -- 78
        44675 => X"4B",  -- 75
        44676 => X"4D",  -- 77
        44677 => X"4A",  -- 74
        44678 => X"47",  -- 71
        44679 => X"4D",  -- 77
        44680 => X"4E",  -- 78
        44681 => X"4F",  -- 79
        44682 => X"4E",  -- 78
        44683 => X"4C",  -- 76
        44684 => X"48",  -- 72
        44685 => X"45",  -- 69
        44686 => X"43",  -- 67
        44687 => X"43",  -- 67
        44688 => X"45",  -- 69
        44689 => X"45",  -- 69
        44690 => X"44",  -- 68
        44691 => X"46",  -- 70
        44692 => X"49",  -- 73
        44693 => X"4B",  -- 75
        44694 => X"48",  -- 72
        44695 => X"44",  -- 68
        44696 => X"43",  -- 67
        44697 => X"43",  -- 67
        44698 => X"40",  -- 64
        44699 => X"3D",  -- 61
        44700 => X"3F",  -- 63
        44701 => X"44",  -- 68
        44702 => X"46",  -- 70
        44703 => X"44",  -- 68
        44704 => X"42",  -- 66
        44705 => X"42",  -- 66
        44706 => X"44",  -- 68
        44707 => X"44",  -- 68
        44708 => X"42",  -- 66
        44709 => X"48",  -- 72
        44710 => X"5A",  -- 90
        44711 => X"6C",  -- 108
        44712 => X"7F",  -- 127
        44713 => X"94",  -- 148
        44714 => X"9E",  -- 158
        44715 => X"9F",  -- 159
        44716 => X"A9",  -- 169
        44717 => X"AA",  -- 170
        44718 => X"9B",  -- 155
        44719 => X"8F",  -- 143
        44720 => X"8F",  -- 143
        44721 => X"8C",  -- 140
        44722 => X"93",  -- 147
        44723 => X"A4",  -- 164
        44724 => X"B0",  -- 176
        44725 => X"AD",  -- 173
        44726 => X"A3",  -- 163
        44727 => X"9E",  -- 158
        44728 => X"AB",  -- 171
        44729 => X"A5",  -- 165
        44730 => X"A4",  -- 164
        44731 => X"98",  -- 152
        44732 => X"A3",  -- 163
        44733 => X"9C",  -- 156
        44734 => X"9A",  -- 154
        44735 => X"8B",  -- 139
        44736 => X"98",  -- 152
        44737 => X"AF",  -- 175
        44738 => X"A2",  -- 162
        44739 => X"A8",  -- 168
        44740 => X"A8",  -- 168
        44741 => X"AF",  -- 175
        44742 => X"A2",  -- 162
        44743 => X"97",  -- 151
        44744 => X"8F",  -- 143
        44745 => X"90",  -- 144
        44746 => X"92",  -- 146
        44747 => X"97",  -- 151
        44748 => X"9E",  -- 158
        44749 => X"A8",  -- 168
        44750 => X"AC",  -- 172
        44751 => X"AC",  -- 172
        44752 => X"B2",  -- 178
        44753 => X"B0",  -- 176
        44754 => X"B0",  -- 176
        44755 => X"B1",  -- 177
        44756 => X"AF",  -- 175
        44757 => X"B1",  -- 177
        44758 => X"B2",  -- 178
        44759 => X"B5",  -- 181
        44760 => X"AC",  -- 172
        44761 => X"A9",  -- 169
        44762 => X"A8",  -- 168
        44763 => X"AF",  -- 175
        44764 => X"B7",  -- 183
        44765 => X"BB",  -- 187
        44766 => X"BB",  -- 187
        44767 => X"BE",  -- 190
        44768 => X"C6",  -- 198
        44769 => X"CA",  -- 202
        44770 => X"C7",  -- 199
        44771 => X"BE",  -- 190
        44772 => X"BE",  -- 190
        44773 => X"C6",  -- 198
        44774 => X"CA",  -- 202
        44775 => X"C8",  -- 200
        44776 => X"C2",  -- 194
        44777 => X"BB",  -- 187
        44778 => X"B3",  -- 179
        44779 => X"AE",  -- 174
        44780 => X"AB",  -- 171
        44781 => X"A5",  -- 165
        44782 => X"98",  -- 152
        44783 => X"8E",  -- 142
        44784 => X"6D",  -- 109
        44785 => X"53",  -- 83
        44786 => X"3D",  -- 61
        44787 => X"2E",  -- 46
        44788 => X"24",  -- 36
        44789 => X"36",  -- 54
        44790 => X"4C",  -- 76
        44791 => X"4C",  -- 76
        44792 => X"55",  -- 85
        44793 => X"78",  -- 120
        44794 => X"91",  -- 145
        44795 => X"94",  -- 148
        44796 => X"95",  -- 149
        44797 => X"82",  -- 130
        44798 => X"5F",  -- 95
        44799 => X"49",  -- 73
        44800 => X"64",  -- 100
        44801 => X"69",  -- 105
        44802 => X"6E",  -- 110
        44803 => X"73",  -- 115
        44804 => X"77",  -- 119
        44805 => X"7B",  -- 123
        44806 => X"7E",  -- 126
        44807 => X"80",  -- 128
        44808 => X"7D",  -- 125
        44809 => X"7B",  -- 123
        44810 => X"78",  -- 120
        44811 => X"75",  -- 117
        44812 => X"73",  -- 115
        44813 => X"70",  -- 112
        44814 => X"6C",  -- 108
        44815 => X"6A",  -- 106
        44816 => X"67",  -- 103
        44817 => X"63",  -- 99
        44818 => X"5E",  -- 94
        44819 => X"57",  -- 87
        44820 => X"51",  -- 81
        44821 => X"4F",  -- 79
        44822 => X"4F",  -- 79
        44823 => X"4E",  -- 78
        44824 => X"58",  -- 88
        44825 => X"5D",  -- 93
        44826 => X"5E",  -- 94
        44827 => X"5E",  -- 94
        44828 => X"5E",  -- 94
        44829 => X"59",  -- 89
        44830 => X"5E",  -- 94
        44831 => X"6F",  -- 111
        44832 => X"6F",  -- 111
        44833 => X"7E",  -- 126
        44834 => X"68",  -- 104
        44835 => X"6F",  -- 111
        44836 => X"56",  -- 86
        44837 => X"49",  -- 73
        44838 => X"41",  -- 65
        44839 => X"34",  -- 52
        44840 => X"31",  -- 49
        44841 => X"38",  -- 56
        44842 => X"57",  -- 87
        44843 => X"4C",  -- 76
        44844 => X"24",  -- 36
        44845 => X"12",  -- 18
        44846 => X"09",  -- 9
        44847 => X"03",  -- 3
        44848 => X"05",  -- 5
        44849 => X"12",  -- 18
        44850 => X"10",  -- 16
        44851 => X"0E",  -- 14
        44852 => X"14",  -- 20
        44853 => X"12",  -- 18
        44854 => X"32",  -- 50
        44855 => X"6D",  -- 109
        44856 => X"4A",  -- 74
        44857 => X"1D",  -- 29
        44858 => X"35",  -- 53
        44859 => X"48",  -- 72
        44860 => X"56",  -- 86
        44861 => X"6A",  -- 106
        44862 => X"5C",  -- 92
        44863 => X"61",  -- 97
        44864 => X"61",  -- 97
        44865 => X"60",  -- 96
        44866 => X"6D",  -- 109
        44867 => X"5D",  -- 93
        44868 => X"4D",  -- 77
        44869 => X"3D",  -- 61
        44870 => X"2A",  -- 42
        44871 => X"3F",  -- 63
        44872 => X"46",  -- 70
        44873 => X"3C",  -- 60
        44874 => X"38",  -- 56
        44875 => X"37",  -- 55
        44876 => X"2E",  -- 46
        44877 => X"23",  -- 35
        44878 => X"28",  -- 40
        44879 => X"39",  -- 57
        44880 => X"46",  -- 70
        44881 => X"44",  -- 68
        44882 => X"48",  -- 72
        44883 => X"58",  -- 88
        44884 => X"67",  -- 103
        44885 => X"6D",  -- 109
        44886 => X"69",  -- 105
        44887 => X"66",  -- 102
        44888 => X"74",  -- 116
        44889 => X"6E",  -- 110
        44890 => X"7B",  -- 123
        44891 => X"7A",  -- 122
        44892 => X"7A",  -- 122
        44893 => X"75",  -- 117
        44894 => X"7F",  -- 127
        44895 => X"76",  -- 118
        44896 => X"6D",  -- 109
        44897 => X"83",  -- 131
        44898 => X"84",  -- 132
        44899 => X"7E",  -- 126
        44900 => X"87",  -- 135
        44901 => X"8B",  -- 139
        44902 => X"82",  -- 130
        44903 => X"97",  -- 151
        44904 => X"82",  -- 130
        44905 => X"91",  -- 145
        44906 => X"7D",  -- 125
        44907 => X"6A",  -- 106
        44908 => X"66",  -- 102
        44909 => X"65",  -- 101
        44910 => X"63",  -- 99
        44911 => X"53",  -- 83
        44912 => X"52",  -- 82
        44913 => X"51",  -- 81
        44914 => X"63",  -- 99
        44915 => X"5A",  -- 90
        44916 => X"51",  -- 81
        44917 => X"4D",  -- 77
        44918 => X"66",  -- 102
        44919 => X"67",  -- 103
        44920 => X"75",  -- 117
        44921 => X"82",  -- 130
        44922 => X"8F",  -- 143
        44923 => X"94",  -- 148
        44924 => X"93",  -- 147
        44925 => X"8F",  -- 143
        44926 => X"85",  -- 133
        44927 => X"7E",  -- 126
        44928 => X"73",  -- 115
        44929 => X"92",  -- 146
        44930 => X"95",  -- 149
        44931 => X"83",  -- 131
        44932 => X"50",  -- 80
        44933 => X"2A",  -- 42
        44934 => X"53",  -- 83
        44935 => X"83",  -- 131
        44936 => X"4B",  -- 75
        44937 => X"45",  -- 69
        44938 => X"55",  -- 85
        44939 => X"21",  -- 33
        44940 => X"19",  -- 25
        44941 => X"1E",  -- 30
        44942 => X"18",  -- 24
        44943 => X"22",  -- 34
        44944 => X"1F",  -- 31
        44945 => X"16",  -- 22
        44946 => X"15",  -- 21
        44947 => X"22",  -- 34
        44948 => X"5F",  -- 95
        44949 => X"88",  -- 136
        44950 => X"A2",  -- 162
        44951 => X"9F",  -- 159
        44952 => X"80",  -- 128
        44953 => X"64",  -- 100
        44954 => X"4E",  -- 78
        44955 => X"4F",  -- 79
        44956 => X"66",  -- 102
        44957 => X"64",  -- 100
        44958 => X"6B",  -- 107
        44959 => X"7D",  -- 125
        44960 => X"83",  -- 131
        44961 => X"8D",  -- 141
        44962 => X"80",  -- 128
        44963 => X"83",  -- 131
        44964 => X"9F",  -- 159
        44965 => X"B0",  -- 176
        44966 => X"AC",  -- 172
        44967 => X"B5",  -- 181
        44968 => X"CC",  -- 204
        44969 => X"CD",  -- 205
        44970 => X"9E",  -- 158
        44971 => X"A8",  -- 168
        44972 => X"C0",  -- 192
        44973 => X"90",  -- 144
        44974 => X"5D",  -- 93
        44975 => X"4C",  -- 76
        44976 => X"49",  -- 73
        44977 => X"48",  -- 72
        44978 => X"46",  -- 70
        44979 => X"45",  -- 69
        44980 => X"46",  -- 70
        44981 => X"46",  -- 70
        44982 => X"46",  -- 70
        44983 => X"46",  -- 70
        44984 => X"40",  -- 64
        44985 => X"43",  -- 67
        44986 => X"49",  -- 73
        44987 => X"4E",  -- 78
        44988 => X"51",  -- 81
        44989 => X"52",  -- 82
        44990 => X"4E",  -- 78
        44991 => X"4D",  -- 77
        44992 => X"48",  -- 72
        44993 => X"4E",  -- 78
        44994 => X"4B",  -- 75
        44995 => X"49",  -- 73
        44996 => X"4C",  -- 76
        44997 => X"49",  -- 73
        44998 => X"46",  -- 70
        44999 => X"4C",  -- 76
        45000 => X"4C",  -- 76
        45001 => X"4D",  -- 77
        45002 => X"4E",  -- 78
        45003 => X"4C",  -- 76
        45004 => X"49",  -- 73
        45005 => X"45",  -- 69
        45006 => X"42",  -- 66
        45007 => X"42",  -- 66
        45008 => X"43",  -- 67
        45009 => X"42",  -- 66
        45010 => X"42",  -- 66
        45011 => X"44",  -- 68
        45012 => X"46",  -- 70
        45013 => X"46",  -- 70
        45014 => X"44",  -- 68
        45015 => X"42",  -- 66
        45016 => X"44",  -- 68
        45017 => X"43",  -- 67
        45018 => X"40",  -- 64
        45019 => X"3C",  -- 60
        45020 => X"3E",  -- 62
        45021 => X"44",  -- 68
        45022 => X"47",  -- 71
        45023 => X"46",  -- 70
        45024 => X"41",  -- 65
        45025 => X"41",  -- 65
        45026 => X"42",  -- 66
        45027 => X"42",  -- 66
        45028 => X"43",  -- 67
        45029 => X"4D",  -- 77
        45030 => X"60",  -- 96
        45031 => X"70",  -- 112
        45032 => X"7E",  -- 126
        45033 => X"92",  -- 146
        45034 => X"9B",  -- 155
        45035 => X"9E",  -- 158
        45036 => X"A9",  -- 169
        45037 => X"AB",  -- 171
        45038 => X"9F",  -- 159
        45039 => X"96",  -- 150
        45040 => X"91",  -- 145
        45041 => X"92",  -- 146
        45042 => X"99",  -- 153
        45043 => X"A5",  -- 165
        45044 => X"AF",  -- 175
        45045 => X"B1",  -- 177
        45046 => X"AA",  -- 170
        45047 => X"A2",  -- 162
        45048 => X"A8",  -- 168
        45049 => X"A5",  -- 165
        45050 => X"A8",  -- 168
        45051 => X"9C",  -- 156
        45052 => X"A5",  -- 165
        45053 => X"9B",  -- 155
        45054 => X"9E",  -- 158
        45055 => X"96",  -- 150
        45056 => X"92",  -- 146
        45057 => X"AF",  -- 175
        45058 => X"A4",  -- 164
        45059 => X"A4",  -- 164
        45060 => X"A1",  -- 161
        45061 => X"B4",  -- 180
        45062 => X"AD",  -- 173
        45063 => X"9A",  -- 154
        45064 => X"9B",  -- 155
        45065 => X"98",  -- 152
        45066 => X"98",  -- 152
        45067 => X"9D",  -- 157
        45068 => X"A3",  -- 163
        45069 => X"A7",  -- 167
        45070 => X"AA",  -- 170
        45071 => X"AA",  -- 170
        45072 => X"B1",  -- 177
        45073 => X"B5",  -- 181
        45074 => X"B5",  -- 181
        45075 => X"B2",  -- 178
        45076 => X"AD",  -- 173
        45077 => X"AE",  -- 174
        45078 => X"B1",  -- 177
        45079 => X"B5",  -- 181
        45080 => X"AB",  -- 171
        45081 => X"A7",  -- 167
        45082 => X"A9",  -- 169
        45083 => X"AF",  -- 175
        45084 => X"B5",  -- 181
        45085 => X"B9",  -- 185
        45086 => X"BD",  -- 189
        45087 => X"C1",  -- 193
        45088 => X"C0",  -- 192
        45089 => X"C9",  -- 201
        45090 => X"CA",  -- 202
        45091 => X"BF",  -- 191
        45092 => X"B8",  -- 184
        45093 => X"BC",  -- 188
        45094 => X"C4",  -- 196
        45095 => X"C8",  -- 200
        45096 => X"C4",  -- 196
        45097 => X"BC",  -- 188
        45098 => X"B3",  -- 179
        45099 => X"AB",  -- 171
        45100 => X"A4",  -- 164
        45101 => X"A1",  -- 161
        45102 => X"A0",  -- 160
        45103 => X"A1",  -- 161
        45104 => X"78",  -- 120
        45105 => X"55",  -- 85
        45106 => X"3C",  -- 60
        45107 => X"2F",  -- 47
        45108 => X"24",  -- 36
        45109 => X"2F",  -- 47
        45110 => X"46",  -- 70
        45111 => X"4D",  -- 77
        45112 => X"60",  -- 96
        45113 => X"6B",  -- 107
        45114 => X"7A",  -- 122
        45115 => X"8B",  -- 139
        45116 => X"97",  -- 151
        45117 => X"8A",  -- 138
        45118 => X"68",  -- 104
        45119 => X"4F",  -- 79
        45120 => X"63",  -- 99
        45121 => X"68",  -- 104
        45122 => X"6E",  -- 110
        45123 => X"71",  -- 113
        45124 => X"74",  -- 116
        45125 => X"78",  -- 120
        45126 => X"7D",  -- 125
        45127 => X"81",  -- 129
        45128 => X"85",  -- 133
        45129 => X"85",  -- 133
        45130 => X"81",  -- 129
        45131 => X"7C",  -- 124
        45132 => X"75",  -- 117
        45133 => X"6E",  -- 110
        45134 => X"68",  -- 104
        45135 => X"66",  -- 102
        45136 => X"67",  -- 103
        45137 => X"62",  -- 98
        45138 => X"5D",  -- 93
        45139 => X"59",  -- 89
        45140 => X"55",  -- 85
        45141 => X"52",  -- 82
        45142 => X"4D",  -- 77
        45143 => X"4B",  -- 75
        45144 => X"50",  -- 80
        45145 => X"54",  -- 84
        45146 => X"52",  -- 82
        45147 => X"54",  -- 84
        45148 => X"59",  -- 89
        45149 => X"58",  -- 88
        45150 => X"5A",  -- 90
        45151 => X"65",  -- 101
        45152 => X"69",  -- 105
        45153 => X"7C",  -- 124
        45154 => X"6A",  -- 106
        45155 => X"75",  -- 117
        45156 => X"59",  -- 89
        45157 => X"61",  -- 97
        45158 => X"4C",  -- 76
        45159 => X"42",  -- 66
        45160 => X"3A",  -- 58
        45161 => X"3A",  -- 58
        45162 => X"5B",  -- 91
        45163 => X"60",  -- 96
        45164 => X"44",  -- 68
        45165 => X"29",  -- 41
        45166 => X"12",  -- 18
        45167 => X"08",  -- 8
        45168 => X"09",  -- 9
        45169 => X"11",  -- 17
        45170 => X"0F",  -- 15
        45171 => X"0F",  -- 15
        45172 => X"12",  -- 18
        45173 => X"0F",  -- 15
        45174 => X"20",  -- 32
        45175 => X"44",  -- 68
        45176 => X"26",  -- 38
        45177 => X"00",  -- 0
        45178 => X"2D",  -- 45
        45179 => X"72",  -- 114
        45180 => X"80",  -- 128
        45181 => X"6F",  -- 111
        45182 => X"58",  -- 88
        45183 => X"5F",  -- 95
        45184 => X"64",  -- 100
        45185 => X"62",  -- 98
        45186 => X"61",  -- 97
        45187 => X"52",  -- 82
        45188 => X"44",  -- 68
        45189 => X"36",  -- 54
        45190 => X"33",  -- 51
        45191 => X"4A",  -- 74
        45192 => X"44",  -- 68
        45193 => X"3C",  -- 60
        45194 => X"37",  -- 55
        45195 => X"34",  -- 52
        45196 => X"2C",  -- 44
        45197 => X"26",  -- 38
        45198 => X"2E",  -- 46
        45199 => X"3E",  -- 62
        45200 => X"48",  -- 72
        45201 => X"4B",  -- 75
        45202 => X"53",  -- 83
        45203 => X"5D",  -- 93
        45204 => X"63",  -- 99
        45205 => X"64",  -- 100
        45206 => X"64",  -- 100
        45207 => X"65",  -- 101
        45208 => X"69",  -- 105
        45209 => X"68",  -- 104
        45210 => X"76",  -- 118
        45211 => X"72",  -- 114
        45212 => X"82",  -- 130
        45213 => X"77",  -- 119
        45214 => X"81",  -- 129
        45215 => X"82",  -- 130
        45216 => X"6C",  -- 108
        45217 => X"89",  -- 137
        45218 => X"7A",  -- 122
        45219 => X"7E",  -- 126
        45220 => X"7E",  -- 126
        45221 => X"83",  -- 131
        45222 => X"8B",  -- 139
        45223 => X"8D",  -- 141
        45224 => X"7E",  -- 126
        45225 => X"8C",  -- 140
        45226 => X"7E",  -- 126
        45227 => X"70",  -- 112
        45228 => X"6C",  -- 108
        45229 => X"67",  -- 103
        45230 => X"68",  -- 104
        45231 => X"61",  -- 97
        45232 => X"59",  -- 89
        45233 => X"69",  -- 105
        45234 => X"65",  -- 101
        45235 => X"52",  -- 82
        45236 => X"5F",  -- 95
        45237 => X"4C",  -- 76
        45238 => X"4E",  -- 78
        45239 => X"69",  -- 105
        45240 => X"7A",  -- 122
        45241 => X"83",  -- 131
        45242 => X"89",  -- 137
        45243 => X"89",  -- 137
        45244 => X"89",  -- 137
        45245 => X"8D",  -- 141
        45246 => X"90",  -- 144
        45247 => X"8E",  -- 142
        45248 => X"91",  -- 145
        45249 => X"86",  -- 134
        45250 => X"97",  -- 151
        45251 => X"89",  -- 137
        45252 => X"5A",  -- 90
        45253 => X"55",  -- 85
        45254 => X"64",  -- 100
        45255 => X"55",  -- 85
        45256 => X"20",  -- 32
        45257 => X"27",  -- 39
        45258 => X"3D",  -- 61
        45259 => X"23",  -- 35
        45260 => X"19",  -- 25
        45261 => X"1D",  -- 29
        45262 => X"15",  -- 21
        45263 => X"1A",  -- 26
        45264 => X"13",  -- 19
        45265 => X"13",  -- 19
        45266 => X"17",  -- 23
        45267 => X"1C",  -- 28
        45268 => X"51",  -- 81
        45269 => X"7F",  -- 127
        45270 => X"91",  -- 145
        45271 => X"7C",  -- 124
        45272 => X"50",  -- 80
        45273 => X"51",  -- 81
        45274 => X"50",  -- 80
        45275 => X"53",  -- 83
        45276 => X"6F",  -- 111
        45277 => X"6E",  -- 110
        45278 => X"76",  -- 118
        45279 => X"86",  -- 134
        45280 => X"8A",  -- 138
        45281 => X"9A",  -- 154
        45282 => X"8D",  -- 141
        45283 => X"7C",  -- 124
        45284 => X"A8",  -- 168
        45285 => X"B1",  -- 177
        45286 => X"AF",  -- 175
        45287 => X"B3",  -- 179
        45288 => X"C7",  -- 199
        45289 => X"D3",  -- 211
        45290 => X"A7",  -- 167
        45291 => X"97",  -- 151
        45292 => X"B1",  -- 177
        45293 => X"90",  -- 144
        45294 => X"5D",  -- 93
        45295 => X"52",  -- 82
        45296 => X"49",  -- 73
        45297 => X"47",  -- 71
        45298 => X"46",  -- 70
        45299 => X"46",  -- 70
        45300 => X"47",  -- 71
        45301 => X"47",  -- 71
        45302 => X"46",  -- 70
        45303 => X"45",  -- 69
        45304 => X"41",  -- 65
        45305 => X"42",  -- 66
        45306 => X"47",  -- 71
        45307 => X"4D",  -- 77
        45308 => X"51",  -- 81
        45309 => X"51",  -- 81
        45310 => X"4C",  -- 76
        45311 => X"48",  -- 72
        45312 => X"45",  -- 69
        45313 => X"4A",  -- 74
        45314 => X"47",  -- 71
        45315 => X"46",  -- 70
        45316 => X"4A",  -- 74
        45317 => X"48",  -- 72
        45318 => X"44",  -- 68
        45319 => X"48",  -- 72
        45320 => X"48",  -- 72
        45321 => X"4A",  -- 74
        45322 => X"4C",  -- 76
        45323 => X"4C",  -- 76
        45324 => X"49",  -- 73
        45325 => X"45",  -- 69
        45326 => X"42",  -- 66
        45327 => X"41",  -- 65
        45328 => X"42",  -- 66
        45329 => X"40",  -- 64
        45330 => X"40",  -- 64
        45331 => X"43",  -- 67
        45332 => X"44",  -- 68
        45333 => X"42",  -- 66
        45334 => X"40",  -- 64
        45335 => X"40",  -- 64
        45336 => X"44",  -- 68
        45337 => X"43",  -- 67
        45338 => X"40",  -- 64
        45339 => X"3C",  -- 60
        45340 => X"3E",  -- 62
        45341 => X"44",  -- 68
        45342 => X"47",  -- 71
        45343 => X"46",  -- 70
        45344 => X"41",  -- 65
        45345 => X"42",  -- 66
        45346 => X"41",  -- 65
        45347 => X"40",  -- 64
        45348 => X"44",  -- 68
        45349 => X"50",  -- 80
        45350 => X"66",  -- 102
        45351 => X"76",  -- 118
        45352 => X"81",  -- 129
        45353 => X"90",  -- 144
        45354 => X"98",  -- 152
        45355 => X"9E",  -- 158
        45356 => X"A8",  -- 168
        45357 => X"A7",  -- 167
        45358 => X"9E",  -- 158
        45359 => X"9A",  -- 154
        45360 => X"94",  -- 148
        45361 => X"93",  -- 147
        45362 => X"98",  -- 152
        45363 => X"A1",  -- 161
        45364 => X"A6",  -- 166
        45365 => X"A6",  -- 166
        45366 => X"A2",  -- 162
        45367 => X"9E",  -- 158
        45368 => X"A1",  -- 161
        45369 => X"A2",  -- 162
        45370 => X"A7",  -- 167
        45371 => X"A0",  -- 160
        45372 => X"A2",  -- 162
        45373 => X"9D",  -- 157
        45374 => X"A0",  -- 160
        45375 => X"9F",  -- 159
        45376 => X"92",  -- 146
        45377 => X"AC",  -- 172
        45378 => X"A2",  -- 162
        45379 => X"A1",  -- 161
        45380 => X"9D",  -- 157
        45381 => X"B2",  -- 178
        45382 => X"B5",  -- 181
        45383 => X"A4",  -- 164
        45384 => X"AD",  -- 173
        45385 => X"A5",  -- 165
        45386 => X"A0",  -- 160
        45387 => X"A2",  -- 162
        45388 => X"A5",  -- 165
        45389 => X"A4",  -- 164
        45390 => X"A8",  -- 168
        45391 => X"AB",  -- 171
        45392 => X"AF",  -- 175
        45393 => X"B5",  -- 181
        45394 => X"B6",  -- 182
        45395 => X"B2",  -- 178
        45396 => X"AC",  -- 172
        45397 => X"A8",  -- 168
        45398 => X"A9",  -- 169
        45399 => X"A9",  -- 169
        45400 => X"AB",  -- 171
        45401 => X"AB",  -- 171
        45402 => X"AD",  -- 173
        45403 => X"B4",  -- 180
        45404 => X"B8",  -- 184
        45405 => X"BA",  -- 186
        45406 => X"BF",  -- 191
        45407 => X"C6",  -- 198
        45408 => X"C1",  -- 193
        45409 => X"C7",  -- 199
        45410 => X"CA",  -- 202
        45411 => X"C4",  -- 196
        45412 => X"BA",  -- 186
        45413 => X"B7",  -- 183
        45414 => X"BD",  -- 189
        45415 => X"C5",  -- 197
        45416 => X"C4",  -- 196
        45417 => X"BF",  -- 191
        45418 => X"B6",  -- 182
        45419 => X"AC",  -- 172
        45420 => X"A0",  -- 160
        45421 => X"9A",  -- 154
        45422 => X"9C",  -- 156
        45423 => X"A3",  -- 163
        45424 => X"A3",  -- 163
        45425 => X"5F",  -- 95
        45426 => X"2D",  -- 45
        45427 => X"2B",  -- 43
        45428 => X"2D",  -- 45
        45429 => X"29",  -- 41
        45430 => X"36",  -- 54
        45431 => X"4A",  -- 74
        45432 => X"54",  -- 84
        45433 => X"5E",  -- 94
        45434 => X"75",  -- 117
        45435 => X"84",  -- 132
        45436 => X"83",  -- 131
        45437 => X"77",  -- 119
        45438 => X"6F",  -- 111
        45439 => X"70",  -- 112
        45440 => X"66",  -- 102
        45441 => X"6A",  -- 106
        45442 => X"71",  -- 113
        45443 => X"72",  -- 114
        45444 => X"72",  -- 114
        45445 => X"73",  -- 115
        45446 => X"76",  -- 118
        45447 => X"7A",  -- 122
        45448 => X"80",  -- 128
        45449 => X"82",  -- 130
        45450 => X"83",  -- 131
        45451 => X"7E",  -- 126
        45452 => X"74",  -- 116
        45453 => X"6C",  -- 108
        45454 => X"68",  -- 104
        45455 => X"68",  -- 104
        45456 => X"67",  -- 103
        45457 => X"64",  -- 100
        45458 => X"5F",  -- 95
        45459 => X"5E",  -- 94
        45460 => X"5D",  -- 93
        45461 => X"5B",  -- 91
        45462 => X"53",  -- 83
        45463 => X"4F",  -- 79
        45464 => X"4A",  -- 74
        45465 => X"4D",  -- 77
        45466 => X"4A",  -- 74
        45467 => X"4A",  -- 74
        45468 => X"50",  -- 80
        45469 => X"52",  -- 82
        45470 => X"55",  -- 85
        45471 => X"60",  -- 96
        45472 => X"6A",  -- 106
        45473 => X"6F",  -- 111
        45474 => X"70",  -- 112
        45475 => X"77",  -- 119
        45476 => X"6A",  -- 106
        45477 => X"6F",  -- 111
        45478 => X"54",  -- 84
        45479 => X"4D",  -- 77
        45480 => X"3C",  -- 60
        45481 => X"3D",  -- 61
        45482 => X"56",  -- 86
        45483 => X"5F",  -- 95
        45484 => X"55",  -- 85
        45485 => X"45",  -- 69
        45486 => X"29",  -- 41
        45487 => X"1D",  -- 29
        45488 => X"10",  -- 16
        45489 => X"0F",  -- 15
        45490 => X"11",  -- 17
        45491 => X"1A",  -- 26
        45492 => X"21",  -- 33
        45493 => X"1F",  -- 31
        45494 => X"1C",  -- 28
        45495 => X"1B",  -- 27
        45496 => X"27",  -- 39
        45497 => X"0C",  -- 12
        45498 => X"3A",  -- 58
        45499 => X"7D",  -- 125
        45500 => X"77",  -- 119
        45501 => X"59",  -- 89
        45502 => X"52",  -- 82
        45503 => X"57",  -- 87
        45504 => X"5E",  -- 94
        45505 => X"5C",  -- 92
        45506 => X"4C",  -- 76
        45507 => X"49",  -- 73
        45508 => X"43",  -- 67
        45509 => X"32",  -- 50
        45510 => X"38",  -- 56
        45511 => X"45",  -- 69
        45512 => X"3D",  -- 61
        45513 => X"3C",  -- 60
        45514 => X"37",  -- 55
        45515 => X"31",  -- 49
        45516 => X"29",  -- 41
        45517 => X"2A",  -- 42
        45518 => X"3B",  -- 59
        45519 => X"4F",  -- 79
        45520 => X"53",  -- 83
        45521 => X"5C",  -- 92
        45522 => X"63",  -- 99
        45523 => X"62",  -- 98
        45524 => X"58",  -- 88
        45525 => X"52",  -- 82
        45526 => X"5C",  -- 92
        45527 => X"69",  -- 105
        45528 => X"5E",  -- 94
        45529 => X"68",  -- 104
        45530 => X"68",  -- 104
        45531 => X"6D",  -- 109
        45532 => X"80",  -- 128
        45533 => X"78",  -- 120
        45534 => X"71",  -- 113
        45535 => X"7C",  -- 124
        45536 => X"6F",  -- 111
        45537 => X"77",  -- 119
        45538 => X"68",  -- 104
        45539 => X"77",  -- 119
        45540 => X"74",  -- 116
        45541 => X"7A",  -- 122
        45542 => X"79",  -- 121
        45543 => X"72",  -- 114
        45544 => X"70",  -- 112
        45545 => X"82",  -- 130
        45546 => X"7E",  -- 126
        45547 => X"78",  -- 120
        45548 => X"72",  -- 114
        45549 => X"67",  -- 103
        45550 => X"6C",  -- 108
        45551 => X"6F",  -- 111
        45552 => X"59",  -- 89
        45553 => X"62",  -- 98
        45554 => X"5F",  -- 95
        45555 => X"56",  -- 86
        45556 => X"6B",  -- 107
        45557 => X"4F",  -- 79
        45558 => X"45",  -- 69
        45559 => X"58",  -- 88
        45560 => X"75",  -- 117
        45561 => X"7D",  -- 125
        45562 => X"80",  -- 128
        45563 => X"7F",  -- 127
        45564 => X"84",  -- 132
        45565 => X"90",  -- 144
        45566 => X"94",  -- 148
        45567 => X"90",  -- 144
        45568 => X"A6",  -- 166
        45569 => X"9F",  -- 159
        45570 => X"95",  -- 149
        45571 => X"68",  -- 104
        45572 => X"67",  -- 103
        45573 => X"7D",  -- 125
        45574 => X"49",  -- 73
        45575 => X"17",  -- 23
        45576 => X"15",  -- 21
        45577 => X"2D",  -- 45
        45578 => X"40",  -- 64
        45579 => X"35",  -- 53
        45580 => X"15",  -- 21
        45581 => X"12",  -- 18
        45582 => X"12",  -- 18
        45583 => X"13",  -- 19
        45584 => X"14",  -- 20
        45585 => X"12",  -- 18
        45586 => X"18",  -- 24
        45587 => X"1E",  -- 30
        45588 => X"4F",  -- 79
        45589 => X"75",  -- 117
        45590 => X"7A",  -- 122
        45591 => X"56",  -- 86
        45592 => X"40",  -- 64
        45593 => X"59",  -- 89
        45594 => X"58",  -- 88
        45595 => X"62",  -- 98
        45596 => X"73",  -- 115
        45597 => X"83",  -- 131
        45598 => X"7D",  -- 125
        45599 => X"8D",  -- 141
        45600 => X"95",  -- 149
        45601 => X"9C",  -- 156
        45602 => X"97",  -- 151
        45603 => X"88",  -- 136
        45604 => X"A2",  -- 162
        45605 => X"AF",  -- 175
        45606 => X"B8",  -- 184
        45607 => X"B8",  -- 184
        45608 => X"BD",  -- 189
        45609 => X"C9",  -- 201
        45610 => X"B9",  -- 185
        45611 => X"94",  -- 148
        45612 => X"91",  -- 145
        45613 => X"88",  -- 136
        45614 => X"62",  -- 98
        45615 => X"52",  -- 82
        45616 => X"4A",  -- 74
        45617 => X"46",  -- 70
        45618 => X"45",  -- 69
        45619 => X"46",  -- 70
        45620 => X"48",  -- 72
        45621 => X"49",  -- 73
        45622 => X"46",  -- 70
        45623 => X"43",  -- 67
        45624 => X"41",  -- 65
        45625 => X"41",  -- 65
        45626 => X"44",  -- 68
        45627 => X"4A",  -- 74
        45628 => X"4E",  -- 78
        45629 => X"4E",  -- 78
        45630 => X"49",  -- 73
        45631 => X"44",  -- 68
        45632 => X"43",  -- 67
        45633 => X"46",  -- 70
        45634 => X"42",  -- 66
        45635 => X"42",  -- 66
        45636 => X"49",  -- 73
        45637 => X"47",  -- 71
        45638 => X"41",  -- 65
        45639 => X"43",  -- 67
        45640 => X"43",  -- 67
        45641 => X"46",  -- 70
        45642 => X"49",  -- 73
        45643 => X"4A",  -- 74
        45644 => X"48",  -- 72
        45645 => X"45",  -- 69
        45646 => X"42",  -- 66
        45647 => X"41",  -- 65
        45648 => X"43",  -- 67
        45649 => X"40",  -- 64
        45650 => X"40",  -- 64
        45651 => X"43",  -- 67
        45652 => X"43",  -- 67
        45653 => X"3F",  -- 63
        45654 => X"3D",  -- 61
        45655 => X"3F",  -- 63
        45656 => X"44",  -- 68
        45657 => X"44",  -- 68
        45658 => X"40",  -- 64
        45659 => X"3C",  -- 60
        45660 => X"3E",  -- 62
        45661 => X"44",  -- 68
        45662 => X"46",  -- 70
        45663 => X"45",  -- 69
        45664 => X"44",  -- 68
        45665 => X"44",  -- 68
        45666 => X"42",  -- 66
        45667 => X"3F",  -- 63
        45668 => X"44",  -- 68
        45669 => X"53",  -- 83
        45670 => X"69",  -- 105
        45671 => X"7A",  -- 122
        45672 => X"86",  -- 134
        45673 => X"90",  -- 144
        45674 => X"96",  -- 150
        45675 => X"A1",  -- 161
        45676 => X"A7",  -- 167
        45677 => X"9E",  -- 158
        45678 => X"94",  -- 148
        45679 => X"95",  -- 149
        45680 => X"9A",  -- 154
        45681 => X"8D",  -- 141
        45682 => X"8A",  -- 138
        45683 => X"98",  -- 152
        45684 => X"9F",  -- 159
        45685 => X"99",  -- 153
        45686 => X"96",  -- 150
        45687 => X"9C",  -- 156
        45688 => X"9C",  -- 156
        45689 => X"A0",  -- 160
        45690 => X"9E",  -- 158
        45691 => X"A1",  -- 161
        45692 => X"99",  -- 153
        45693 => X"9C",  -- 156
        45694 => X"99",  -- 153
        45695 => X"9D",  -- 157
        45696 => X"99",  -- 153
        45697 => X"A6",  -- 166
        45698 => X"9D",  -- 157
        45699 => X"A3",  -- 163
        45700 => X"9A",  -- 154
        45701 => X"AA",  -- 170
        45702 => X"B7",  -- 183
        45703 => X"B3",  -- 179
        45704 => X"B7",  -- 183
        45705 => X"AE",  -- 174
        45706 => X"A8",  -- 168
        45707 => X"AB",  -- 171
        45708 => X"AA",  -- 170
        45709 => X"A4",  -- 164
        45710 => X"A4",  -- 164
        45711 => X"AB",  -- 171
        45712 => X"AE",  -- 174
        45713 => X"B2",  -- 178
        45714 => X"B0",  -- 176
        45715 => X"AA",  -- 170
        45716 => X"A7",  -- 167
        45717 => X"A6",  -- 166
        45718 => X"A5",  -- 165
        45719 => X"A3",  -- 163
        45720 => X"A5",  -- 165
        45721 => X"AB",  -- 171
        45722 => X"B4",  -- 180
        45723 => X"B9",  -- 185
        45724 => X"BA",  -- 186
        45725 => X"B9",  -- 185
        45726 => X"BE",  -- 190
        45727 => X"C7",  -- 199
        45728 => X"C7",  -- 199
        45729 => X"C6",  -- 198
        45730 => X"C8",  -- 200
        45731 => X"C9",  -- 201
        45732 => X"C1",  -- 193
        45733 => X"B7",  -- 183
        45734 => X"B7",  -- 183
        45735 => X"BF",  -- 191
        45736 => X"C1",  -- 193
        45737 => X"BE",  -- 190
        45738 => X"BA",  -- 186
        45739 => X"B0",  -- 176
        45740 => X"9F",  -- 159
        45741 => X"90",  -- 144
        45742 => X"8A",  -- 138
        45743 => X"8D",  -- 141
        45744 => X"A2",  -- 162
        45745 => X"8C",  -- 140
        45746 => X"53",  -- 83
        45747 => X"21",  -- 33
        45748 => X"1F",  -- 31
        45749 => X"38",  -- 56
        45750 => X"40",  -- 64
        45751 => X"38",  -- 56
        45752 => X"48",  -- 72
        45753 => X"55",  -- 85
        45754 => X"6D",  -- 109
        45755 => X"75",  -- 117
        45756 => X"6A",  -- 106
        45757 => X"66",  -- 102
        45758 => X"73",  -- 115
        45759 => X"82",  -- 130
        45760 => X"66",  -- 102
        45761 => X"6E",  -- 110
        45762 => X"76",  -- 118
        45763 => X"78",  -- 120
        45764 => X"76",  -- 118
        45765 => X"72",  -- 114
        45766 => X"70",  -- 112
        45767 => X"71",  -- 113
        45768 => X"71",  -- 113
        45769 => X"77",  -- 119
        45770 => X"7C",  -- 124
        45771 => X"7A",  -- 122
        45772 => X"72",  -- 114
        45773 => X"6C",  -- 108
        45774 => X"6B",  -- 107
        45775 => X"6D",  -- 109
        45776 => X"67",  -- 103
        45777 => X"63",  -- 99
        45778 => X"61",  -- 97
        45779 => X"63",  -- 99
        45780 => X"65",  -- 101
        45781 => X"63",  -- 99
        45782 => X"5D",  -- 93
        45783 => X"56",  -- 86
        45784 => X"4B",  -- 75
        45785 => X"4D",  -- 77
        45786 => X"49",  -- 73
        45787 => X"45",  -- 69
        45788 => X"49",  -- 73
        45789 => X"4C",  -- 76
        45790 => X"51",  -- 81
        45791 => X"5E",  -- 94
        45792 => X"6D",  -- 109
        45793 => X"63",  -- 99
        45794 => X"75",  -- 117
        45795 => X"78",  -- 120
        45796 => X"79",  -- 121
        45797 => X"73",  -- 115
        45798 => X"55",  -- 85
        45799 => X"56",  -- 86
        45800 => X"44",  -- 68
        45801 => X"44",  -- 68
        45802 => X"50",  -- 80
        45803 => X"52",  -- 82
        45804 => X"56",  -- 86
        45805 => X"55",  -- 85
        45806 => X"3B",  -- 59
        45807 => X"2C",  -- 44
        45808 => X"32",  -- 50
        45809 => X"2E",  -- 46
        45810 => X"37",  -- 55
        45811 => X"43",  -- 67
        45812 => X"48",  -- 72
        45813 => X"47",  -- 71
        45814 => X"37",  -- 55
        45815 => X"21",  -- 33
        45816 => X"36",  -- 54
        45817 => X"2C",  -- 44
        45818 => X"46",  -- 70
        45819 => X"61",  -- 97
        45820 => X"45",  -- 69
        45821 => X"35",  -- 53
        45822 => X"4B",  -- 75
        45823 => X"4A",  -- 74
        45824 => X"57",  -- 87
        45825 => X"55",  -- 85
        45826 => X"40",  -- 64
        45827 => X"49",  -- 73
        45828 => X"49",  -- 73
        45829 => X"33",  -- 51
        45830 => X"3A",  -- 58
        45831 => X"3C",  -- 60
        45832 => X"3A",  -- 58
        45833 => X"3D",  -- 61
        45834 => X"3A",  -- 58
        45835 => X"2E",  -- 46
        45836 => X"26",  -- 38
        45837 => X"2D",  -- 45
        45838 => X"47",  -- 71
        45839 => X"5C",  -- 92
        45840 => X"66",  -- 102
        45841 => X"61",  -- 97
        45842 => X"5B",  -- 91
        45843 => X"56",  -- 86
        45844 => X"52",  -- 82
        45845 => X"4E",  -- 78
        45846 => X"54",  -- 84
        45847 => X"5B",  -- 91
        45848 => X"60",  -- 96
        45849 => X"71",  -- 113
        45850 => X"61",  -- 97
        45851 => X"6D",  -- 109
        45852 => X"7D",  -- 125
        45853 => X"7C",  -- 124
        45854 => X"5E",  -- 94
        45855 => X"6F",  -- 111
        45856 => X"7A",  -- 122
        45857 => X"7E",  -- 126
        45858 => X"81",  -- 129
        45859 => X"91",  -- 145
        45860 => X"7D",  -- 125
        45861 => X"7E",  -- 126
        45862 => X"78",  -- 120
        45863 => X"80",  -- 128
        45864 => X"77",  -- 119
        45865 => X"7D",  -- 125
        45866 => X"71",  -- 113
        45867 => X"77",  -- 119
        45868 => X"7C",  -- 124
        45869 => X"70",  -- 112
        45870 => X"6A",  -- 106
        45871 => X"61",  -- 97
        45872 => X"56",  -- 86
        45873 => X"45",  -- 69
        45874 => X"57",  -- 87
        45875 => X"66",  -- 102
        45876 => X"68",  -- 104
        45877 => X"52",  -- 82
        45878 => X"4F",  -- 79
        45879 => X"43",  -- 67
        45880 => X"64",  -- 100
        45881 => X"6F",  -- 111
        45882 => X"79",  -- 121
        45883 => X"82",  -- 130
        45884 => X"8E",  -- 142
        45885 => X"9A",  -- 154
        45886 => X"98",  -- 152
        45887 => X"8E",  -- 142
        45888 => X"81",  -- 129
        45889 => X"BB",  -- 187
        45890 => X"A0",  -- 160
        45891 => X"46",  -- 70
        45892 => X"70",  -- 112
        45893 => X"86",  -- 134
        45894 => X"28",  -- 40
        45895 => X"18",  -- 24
        45896 => X"20",  -- 32
        45897 => X"48",  -- 72
        45898 => X"5D",  -- 93
        45899 => X"5F",  -- 95
        45900 => X"28",  -- 40
        45901 => X"19",  -- 25
        45902 => X"1B",  -- 27
        45903 => X"17",  -- 23
        45904 => X"18",  -- 24
        45905 => X"11",  -- 17
        45906 => X"17",  -- 23
        45907 => X"21",  -- 33
        45908 => X"4F",  -- 79
        45909 => X"6E",  -- 110
        45910 => X"69",  -- 105
        45911 => X"3B",  -- 59
        45912 => X"3D",  -- 61
        45913 => X"63",  -- 99
        45914 => X"5A",  -- 90
        45915 => X"6D",  -- 109
        45916 => X"75",  -- 117
        45917 => X"97",  -- 151
        45918 => X"86",  -- 134
        45919 => X"96",  -- 150
        45920 => X"9F",  -- 159
        45921 => X"9A",  -- 154
        45922 => X"9A",  -- 154
        45923 => X"99",  -- 153
        45924 => X"98",  -- 152
        45925 => X"AC",  -- 172
        45926 => X"BF",  -- 191
        45927 => X"BD",  -- 189
        45928 => X"BD",  -- 189
        45929 => X"C4",  -- 196
        45930 => X"CC",  -- 204
        45931 => X"9B",  -- 155
        45932 => X"75",  -- 117
        45933 => X"7C",  -- 124
        45934 => X"63",  -- 99
        45935 => X"47",  -- 71
        45936 => X"49",  -- 73
        45937 => X"47",  -- 71
        45938 => X"44",  -- 68
        45939 => X"44",  -- 68
        45940 => X"48",  -- 72
        45941 => X"4A",  -- 74
        45942 => X"46",  -- 70
        45943 => X"42",  -- 66
        45944 => X"41",  -- 65
        45945 => X"40",  -- 64
        45946 => X"42",  -- 66
        45947 => X"48",  -- 72
        45948 => X"4D",  -- 77
        45949 => X"4E",  -- 78
        45950 => X"48",  -- 72
        45951 => X"42",  -- 66
        45952 => X"43",  -- 67
        45953 => X"44",  -- 68
        45954 => X"3F",  -- 63
        45955 => X"3F",  -- 63
        45956 => X"47",  -- 71
        45957 => X"46",  -- 70
        45958 => X"3F",  -- 63
        45959 => X"3F",  -- 63
        45960 => X"40",  -- 64
        45961 => X"43",  -- 67
        45962 => X"47",  -- 71
        45963 => X"49",  -- 73
        45964 => X"47",  -- 71
        45965 => X"44",  -- 68
        45966 => X"41",  -- 65
        45967 => X"40",  -- 64
        45968 => X"43",  -- 67
        45969 => X"40",  -- 64
        45970 => X"40",  -- 64
        45971 => X"43",  -- 67
        45972 => X"43",  -- 67
        45973 => X"3E",  -- 62
        45974 => X"3C",  -- 60
        45975 => X"3E",  -- 62
        45976 => X"44",  -- 68
        45977 => X"44",  -- 68
        45978 => X"41",  -- 65
        45979 => X"3D",  -- 61
        45980 => X"3F",  -- 63
        45981 => X"44",  -- 68
        45982 => X"47",  -- 71
        45983 => X"44",  -- 68
        45984 => X"47",  -- 71
        45985 => X"47",  -- 71
        45986 => X"44",  -- 68
        45987 => X"40",  -- 64
        45988 => X"43",  -- 67
        45989 => X"54",  -- 84
        45990 => X"6B",  -- 107
        45991 => X"7B",  -- 123
        45992 => X"8A",  -- 138
        45993 => X"91",  -- 145
        45994 => X"98",  -- 152
        45995 => X"A2",  -- 162
        45996 => X"A6",  -- 166
        45997 => X"97",  -- 151
        45998 => X"8B",  -- 139
        45999 => X"90",  -- 144
        46000 => X"A1",  -- 161
        46001 => X"86",  -- 134
        46002 => X"81",  -- 129
        46003 => X"98",  -- 152
        46004 => X"A2",  -- 162
        46005 => X"96",  -- 150
        46006 => X"93",  -- 147
        46007 => X"A2",  -- 162
        46008 => X"A0",  -- 160
        46009 => X"A2",  -- 162
        46010 => X"9A",  -- 154
        46011 => X"A4",  -- 164
        46012 => X"96",  -- 150
        46013 => X"9B",  -- 155
        46014 => X"93",  -- 147
        46015 => X"98",  -- 152
        46016 => X"9C",  -- 156
        46017 => X"9C",  -- 156
        46018 => X"93",  -- 147
        46019 => X"A3",  -- 163
        46020 => X"96",  -- 150
        46021 => X"A1",  -- 161
        46022 => X"B2",  -- 178
        46023 => X"BC",  -- 188
        46024 => X"B5",  -- 181
        46025 => X"AF",  -- 175
        46026 => X"AF",  -- 175
        46027 => X"B5",  -- 181
        46028 => X"B0",  -- 176
        46029 => X"A6",  -- 166
        46030 => X"A2",  -- 162
        46031 => X"A7",  -- 167
        46032 => X"B3",  -- 179
        46033 => X"B0",  -- 176
        46034 => X"A7",  -- 167
        46035 => X"A0",  -- 160
        46036 => X"A1",  -- 161
        46037 => X"A7",  -- 167
        46038 => X"A9",  -- 169
        46039 => X"A6",  -- 166
        46040 => X"A0",  -- 160
        46041 => X"A9",  -- 169
        46042 => X"B6",  -- 182
        46043 => X"BC",  -- 188
        46044 => X"BA",  -- 186
        46045 => X"B8",  -- 184
        46046 => X"BD",  -- 189
        46047 => X"C4",  -- 196
        46048 => X"CC",  -- 204
        46049 => X"C5",  -- 197
        46050 => X"C5",  -- 197
        46051 => X"CC",  -- 204
        46052 => X"C8",  -- 200
        46053 => X"BA",  -- 186
        46054 => X"B4",  -- 180
        46055 => X"BA",  -- 186
        46056 => X"BD",  -- 189
        46057 => X"BC",  -- 188
        46058 => X"BA",  -- 186
        46059 => X"B3",  -- 179
        46060 => X"A0",  -- 160
        46061 => X"87",  -- 135
        46062 => X"77",  -- 119
        46063 => X"73",  -- 115
        46064 => X"8B",  -- 139
        46065 => X"99",  -- 153
        46066 => X"81",  -- 129
        46067 => X"4F",  -- 79
        46068 => X"2D",  -- 45
        46069 => X"21",  -- 33
        46070 => X"2E",  -- 46
        46071 => X"4A",  -- 74
        46072 => X"58",  -- 88
        46073 => X"53",  -- 83
        46074 => X"58",  -- 88
        46075 => X"5E",  -- 94
        46076 => X"60",  -- 96
        46077 => X"6B",  -- 107
        46078 => X"71",  -- 113
        46079 => X"6D",  -- 109
        46080 => X"6B",  -- 107
        46081 => X"71",  -- 113
        46082 => X"76",  -- 118
        46083 => X"78",  -- 120
        46084 => X"7B",  -- 123
        46085 => X"7F",  -- 127
        46086 => X"7E",  -- 126
        46087 => X"7A",  -- 122
        46088 => X"72",  -- 114
        46089 => X"71",  -- 113
        46090 => X"73",  -- 115
        46091 => X"79",  -- 121
        46092 => X"7A",  -- 122
        46093 => X"76",  -- 118
        46094 => X"74",  -- 116
        46095 => X"76",  -- 118
        46096 => X"6D",  -- 109
        46097 => X"68",  -- 104
        46098 => X"62",  -- 98
        46099 => X"60",  -- 96
        46100 => X"61",  -- 97
        46101 => X"60",  -- 96
        46102 => X"5F",  -- 95
        46103 => X"5B",  -- 91
        46104 => X"52",  -- 82
        46105 => X"52",  -- 82
        46106 => X"52",  -- 82
        46107 => X"4F",  -- 79
        46108 => X"4C",  -- 76
        46109 => X"4F",  -- 79
        46110 => X"57",  -- 87
        46111 => X"5C",  -- 92
        46112 => X"5D",  -- 93
        46113 => X"68",  -- 104
        46114 => X"70",  -- 112
        46115 => X"78",  -- 120
        46116 => X"7C",  -- 124
        46117 => X"6D",  -- 109
        46118 => X"5D",  -- 93
        46119 => X"5C",  -- 92
        46120 => X"51",  -- 81
        46121 => X"4C",  -- 76
        46122 => X"4D",  -- 77
        46123 => X"52",  -- 82
        46124 => X"58",  -- 88
        46125 => X"4C",  -- 76
        46126 => X"31",  -- 49
        46127 => X"2C",  -- 44
        46128 => X"3A",  -- 58
        46129 => X"44",  -- 68
        46130 => X"52",  -- 82
        46131 => X"5E",  -- 94
        46132 => X"64",  -- 100
        46133 => X"66",  -- 102
        46134 => X"51",  -- 81
        46135 => X"2F",  -- 47
        46136 => X"45",  -- 69
        46137 => X"33",  -- 51
        46138 => X"53",  -- 83
        46139 => X"35",  -- 53
        46140 => X"1D",  -- 29
        46141 => X"4A",  -- 74
        46142 => X"56",  -- 86
        46143 => X"61",  -- 97
        46144 => X"61",  -- 97
        46145 => X"3D",  -- 61
        46146 => X"4C",  -- 76
        46147 => X"64",  -- 100
        46148 => X"4A",  -- 74
        46149 => X"3A",  -- 58
        46150 => X"42",  -- 66
        46151 => X"3B",  -- 59
        46152 => X"34",  -- 52
        46153 => X"3D",  -- 61
        46154 => X"41",  -- 65
        46155 => X"37",  -- 55
        46156 => X"2F",  -- 47
        46157 => X"38",  -- 56
        46158 => X"4A",  -- 74
        46159 => X"57",  -- 87
        46160 => X"53",  -- 83
        46161 => X"4F",  -- 79
        46162 => X"4D",  -- 77
        46163 => X"51",  -- 81
        46164 => X"57",  -- 87
        46165 => X"5C",  -- 92
        46166 => X"5D",  -- 93
        46167 => X"5C",  -- 92
        46168 => X"6B",  -- 107
        46169 => X"71",  -- 113
        46170 => X"72",  -- 114
        46171 => X"6C",  -- 108
        46172 => X"6C",  -- 108
        46173 => X"72",  -- 114
        46174 => X"74",  -- 116
        46175 => X"73",  -- 115
        46176 => X"7A",  -- 122
        46177 => X"80",  -- 128
        46178 => X"7C",  -- 124
        46179 => X"77",  -- 119
        46180 => X"7C",  -- 124
        46181 => X"7D",  -- 125
        46182 => X"79",  -- 121
        46183 => X"7C",  -- 124
        46184 => X"7A",  -- 122
        46185 => X"7F",  -- 127
        46186 => X"7D",  -- 125
        46187 => X"76",  -- 118
        46188 => X"6D",  -- 109
        46189 => X"68",  -- 104
        46190 => X"61",  -- 97
        46191 => X"5A",  -- 90
        46192 => X"4F",  -- 79
        46193 => X"5C",  -- 92
        46194 => X"5B",  -- 91
        46195 => X"55",  -- 85
        46196 => X"5B",  -- 91
        46197 => X"62",  -- 98
        46198 => X"5F",  -- 95
        46199 => X"5B",  -- 91
        46200 => X"65",  -- 101
        46201 => X"76",  -- 118
        46202 => X"75",  -- 117
        46203 => X"86",  -- 134
        46204 => X"8C",  -- 140
        46205 => X"8C",  -- 140
        46206 => X"A0",  -- 160
        46207 => X"9E",  -- 158
        46208 => X"6A",  -- 106
        46209 => X"8C",  -- 140
        46210 => X"9C",  -- 156
        46211 => X"41",  -- 65
        46212 => X"52",  -- 82
        46213 => X"4C",  -- 76
        46214 => X"25",  -- 37
        46215 => X"1C",  -- 28
        46216 => X"37",  -- 55
        46217 => X"72",  -- 114
        46218 => X"7E",  -- 126
        46219 => X"75",  -- 117
        46220 => X"54",  -- 84
        46221 => X"32",  -- 50
        46222 => X"2E",  -- 46
        46223 => X"0C",  -- 12
        46224 => X"09",  -- 9
        46225 => X"18",  -- 24
        46226 => X"0F",  -- 15
        46227 => X"4B",  -- 75
        46228 => X"6B",  -- 107
        46229 => X"4E",  -- 78
        46230 => X"4D",  -- 77
        46231 => X"35",  -- 53
        46232 => X"40",  -- 64
        46233 => X"6D",  -- 109
        46234 => X"5E",  -- 94
        46235 => X"6E",  -- 110
        46236 => X"87",  -- 135
        46237 => X"90",  -- 144
        46238 => X"85",  -- 133
        46239 => X"99",  -- 153
        46240 => X"98",  -- 152
        46241 => X"A2",  -- 162
        46242 => X"A4",  -- 164
        46243 => X"A8",  -- 168
        46244 => X"A3",  -- 163
        46245 => X"AA",  -- 170
        46246 => X"C2",  -- 194
        46247 => X"BF",  -- 191
        46248 => X"CC",  -- 204
        46249 => X"B8",  -- 184
        46250 => X"C5",  -- 197
        46251 => X"A6",  -- 166
        46252 => X"76",  -- 118
        46253 => X"5A",  -- 90
        46254 => X"64",  -- 100
        46255 => X"47",  -- 71
        46256 => X"49",  -- 73
        46257 => X"48",  -- 72
        46258 => X"46",  -- 70
        46259 => X"46",  -- 70
        46260 => X"47",  -- 71
        46261 => X"46",  -- 70
        46262 => X"45",  -- 69
        46263 => X"45",  -- 69
        46264 => X"41",  -- 65
        46265 => X"41",  -- 65
        46266 => X"45",  -- 69
        46267 => X"49",  -- 73
        46268 => X"4A",  -- 74
        46269 => X"47",  -- 71
        46270 => X"47",  -- 71
        46271 => X"4A",  -- 74
        46272 => X"3D",  -- 61
        46273 => X"3E",  -- 62
        46274 => X"3D",  -- 61
        46275 => X"3C",  -- 60
        46276 => X"3F",  -- 63
        46277 => X"43",  -- 67
        46278 => X"3F",  -- 63
        46279 => X"37",  -- 55
        46280 => X"3A",  -- 58
        46281 => X"43",  -- 67
        46282 => X"46",  -- 70
        46283 => X"40",  -- 64
        46284 => X"3F",  -- 63
        46285 => X"45",  -- 69
        46286 => X"46",  -- 70
        46287 => X"43",  -- 67
        46288 => X"40",  -- 64
        46289 => X"3F",  -- 63
        46290 => X"40",  -- 64
        46291 => X"44",  -- 68
        46292 => X"42",  -- 66
        46293 => X"3D",  -- 61
        46294 => X"3B",  -- 59
        46295 => X"3E",  -- 62
        46296 => X"3C",  -- 60
        46297 => X"45",  -- 69
        46298 => X"49",  -- 73
        46299 => X"42",  -- 66
        46300 => X"3D",  -- 61
        46301 => X"41",  -- 65
        46302 => X"45",  -- 69
        46303 => X"45",  -- 69
        46304 => X"44",  -- 68
        46305 => X"4D",  -- 77
        46306 => X"47",  -- 71
        46307 => X"3C",  -- 60
        46308 => X"49",  -- 73
        46309 => X"60",  -- 96
        46310 => X"73",  -- 115
        46311 => X"82",  -- 130
        46312 => X"89",  -- 137
        46313 => X"8C",  -- 140
        46314 => X"94",  -- 148
        46315 => X"91",  -- 145
        46316 => X"98",  -- 152
        46317 => X"9E",  -- 158
        46318 => X"98",  -- 152
        46319 => X"A3",  -- 163
        46320 => X"9A",  -- 154
        46321 => X"80",  -- 128
        46322 => X"77",  -- 119
        46323 => X"91",  -- 145
        46324 => X"A1",  -- 161
        46325 => X"92",  -- 146
        46326 => X"8C",  -- 140
        46327 => X"A0",  -- 160
        46328 => X"A8",  -- 168
        46329 => X"AA",  -- 170
        46330 => X"A1",  -- 161
        46331 => X"A8",  -- 168
        46332 => X"A7",  -- 167
        46333 => X"91",  -- 145
        46334 => X"8E",  -- 142
        46335 => X"94",  -- 148
        46336 => X"9B",  -- 155
        46337 => X"90",  -- 144
        46338 => X"A7",  -- 167
        46339 => X"A2",  -- 162
        46340 => X"8F",  -- 143
        46341 => X"9B",  -- 155
        46342 => X"A8",  -- 168
        46343 => X"BE",  -- 190
        46344 => X"B9",  -- 185
        46345 => X"B1",  -- 177
        46346 => X"B4",  -- 180
        46347 => X"B3",  -- 179
        46348 => X"B6",  -- 182
        46349 => X"B6",  -- 182
        46350 => X"A9",  -- 169
        46351 => X"A9",  -- 169
        46352 => X"AA",  -- 170
        46353 => X"B1",  -- 177
        46354 => X"AC",  -- 172
        46355 => X"A3",  -- 163
        46356 => X"A9",  -- 169
        46357 => X"B6",  -- 182
        46358 => X"B3",  -- 179
        46359 => X"A4",  -- 164
        46360 => X"AA",  -- 170
        46361 => X"B0",  -- 176
        46362 => X"B7",  -- 183
        46363 => X"BB",  -- 187
        46364 => X"BC",  -- 188
        46365 => X"BD",  -- 189
        46366 => X"BE",  -- 190
        46367 => X"C0",  -- 192
        46368 => X"CB",  -- 203
        46369 => X"CB",  -- 203
        46370 => X"CB",  -- 203
        46371 => X"CA",  -- 202
        46372 => X"C7",  -- 199
        46373 => X"C1",  -- 193
        46374 => X"B9",  -- 185
        46375 => X"B4",  -- 180
        46376 => X"BC",  -- 188
        46377 => X"BE",  -- 190
        46378 => X"B8",  -- 184
        46379 => X"AE",  -- 174
        46380 => X"AA",  -- 170
        46381 => X"A0",  -- 160
        46382 => X"7F",  -- 127
        46383 => X"5C",  -- 92
        46384 => X"5F",  -- 95
        46385 => X"7C",  -- 124
        46386 => X"79",  -- 121
        46387 => X"6E",  -- 110
        46388 => X"4D",  -- 77
        46389 => X"2E",  -- 46
        46390 => X"38",  -- 56
        46391 => X"35",  -- 53
        46392 => X"4C",  -- 76
        46393 => X"5C",  -- 92
        46394 => X"69",  -- 105
        46395 => X"6B",  -- 107
        46396 => X"65",  -- 101
        46397 => X"5B",  -- 91
        46398 => X"63",  -- 99
        46399 => X"79",  -- 121
        46400 => X"67",  -- 103
        46401 => X"6C",  -- 108
        46402 => X"6F",  -- 111
        46403 => X"6F",  -- 111
        46404 => X"74",  -- 116
        46405 => X"7C",  -- 124
        46406 => X"82",  -- 130
        46407 => X"83",  -- 131
        46408 => X"7D",  -- 125
        46409 => X"7E",  -- 126
        46410 => X"82",  -- 130
        46411 => X"86",  -- 134
        46412 => X"84",  -- 132
        46413 => X"7D",  -- 125
        46414 => X"7A",  -- 122
        46415 => X"7B",  -- 123
        46416 => X"79",  -- 121
        46417 => X"72",  -- 114
        46418 => X"68",  -- 104
        46419 => X"62",  -- 98
        46420 => X"5F",  -- 95
        46421 => X"5D",  -- 93
        46422 => X"59",  -- 89
        46423 => X"56",  -- 86
        46424 => X"57",  -- 87
        46425 => X"58",  -- 88
        46426 => X"59",  -- 89
        46427 => X"57",  -- 87
        46428 => X"54",  -- 84
        46429 => X"56",  -- 86
        46430 => X"5C",  -- 92
        46431 => X"61",  -- 97
        46432 => X"61",  -- 97
        46433 => X"67",  -- 103
        46434 => X"6D",  -- 109
        46435 => X"78",  -- 120
        46436 => X"7C",  -- 124
        46437 => X"6C",  -- 108
        46438 => X"5F",  -- 95
        46439 => X"60",  -- 96
        46440 => X"5A",  -- 90
        46441 => X"50",  -- 80
        46442 => X"4F",  -- 79
        46443 => X"5A",  -- 90
        46444 => X"66",  -- 102
        46445 => X"54",  -- 84
        46446 => X"29",  -- 41
        46447 => X"0F",  -- 15
        46448 => X"16",  -- 22
        46449 => X"26",  -- 38
        46450 => X"42",  -- 66
        46451 => X"56",  -- 86
        46452 => X"60",  -- 96
        46453 => X"68",  -- 104
        46454 => X"5A",  -- 90
        46455 => X"3E",  -- 62
        46456 => X"1F",  -- 31
        46457 => X"5F",  -- 95
        46458 => X"6B",  -- 107
        46459 => X"24",  -- 36
        46460 => X"3C",  -- 60
        46461 => X"67",  -- 103
        46462 => X"79",  -- 121
        46463 => X"77",  -- 119
        46464 => X"58",  -- 88
        46465 => X"58",  -- 88
        46466 => X"5B",  -- 91
        46467 => X"5B",  -- 91
        46468 => X"4E",  -- 78
        46469 => X"41",  -- 65
        46470 => X"3E",  -- 62
        46471 => X"42",  -- 66
        46472 => X"31",  -- 49
        46473 => X"38",  -- 56
        46474 => X"3A",  -- 58
        46475 => X"35",  -- 53
        46476 => X"30",  -- 48
        46477 => X"3A",  -- 58
        46478 => X"4B",  -- 75
        46479 => X"57",  -- 87
        46480 => X"5C",  -- 92
        46481 => X"79",  -- 121
        46482 => X"69",  -- 105
        46483 => X"59",  -- 89
        46484 => X"6C",  -- 108
        46485 => X"63",  -- 99
        46486 => X"58",  -- 88
        46487 => X"76",  -- 118
        46488 => X"64",  -- 100
        46489 => X"6E",  -- 110
        46490 => X"75",  -- 117
        46491 => X"76",  -- 118
        46492 => X"79",  -- 121
        46493 => X"7C",  -- 124
        46494 => X"78",  -- 120
        46495 => X"71",  -- 113
        46496 => X"69",  -- 105
        46497 => X"73",  -- 115
        46498 => X"74",  -- 116
        46499 => X"73",  -- 115
        46500 => X"79",  -- 121
        46501 => X"76",  -- 118
        46502 => X"6C",  -- 108
        46503 => X"6B",  -- 107
        46504 => X"76",  -- 118
        46505 => X"7C",  -- 124
        46506 => X"7E",  -- 126
        46507 => X"79",  -- 121
        46508 => X"74",  -- 116
        46509 => X"72",  -- 114
        46510 => X"72",  -- 114
        46511 => X"71",  -- 113
        46512 => X"54",  -- 84
        46513 => X"63",  -- 99
        46514 => X"63",  -- 99
        46515 => X"59",  -- 89
        46516 => X"59",  -- 89
        46517 => X"5C",  -- 92
        46518 => X"5E",  -- 94
        46519 => X"64",  -- 100
        46520 => X"67",  -- 103
        46521 => X"79",  -- 121
        46522 => X"7C",  -- 124
        46523 => X"75",  -- 117
        46524 => X"5F",  -- 95
        46525 => X"54",  -- 84
        46526 => X"71",  -- 113
        46527 => X"8E",  -- 142
        46528 => X"7A",  -- 122
        46529 => X"88",  -- 136
        46530 => X"BB",  -- 187
        46531 => X"59",  -- 89
        46532 => X"51",  -- 81
        46533 => X"54",  -- 84
        46534 => X"1C",  -- 28
        46535 => X"2A",  -- 42
        46536 => X"74",  -- 116
        46537 => X"8F",  -- 143
        46538 => X"85",  -- 133
        46539 => X"76",  -- 118
        46540 => X"4B",  -- 75
        46541 => X"22",  -- 34
        46542 => X"2B",  -- 43
        46543 => X"25",  -- 37
        46544 => X"11",  -- 17
        46545 => X"0F",  -- 15
        46546 => X"24",  -- 36
        46547 => X"50",  -- 80
        46548 => X"60",  -- 96
        46549 => X"43",  -- 67
        46550 => X"35",  -- 53
        46551 => X"43",  -- 67
        46552 => X"4D",  -- 77
        46553 => X"71",  -- 113
        46554 => X"68",  -- 104
        46555 => X"70",  -- 112
        46556 => X"84",  -- 132
        46557 => X"85",  -- 133
        46558 => X"82",  -- 130
        46559 => X"92",  -- 146
        46560 => X"9E",  -- 158
        46561 => X"A7",  -- 167
        46562 => X"A9",  -- 169
        46563 => X"AD",  -- 173
        46564 => X"A8",  -- 168
        46565 => X"AE",  -- 174
        46566 => X"C4",  -- 196
        46567 => X"C1",  -- 193
        46568 => X"C7",  -- 199
        46569 => X"B6",  -- 182
        46570 => X"B9",  -- 185
        46571 => X"AD",  -- 173
        46572 => X"86",  -- 134
        46573 => X"57",  -- 87
        46574 => X"4E",  -- 78
        46575 => X"50",  -- 80
        46576 => X"4A",  -- 74
        46577 => X"47",  -- 71
        46578 => X"45",  -- 69
        46579 => X"44",  -- 68
        46580 => X"45",  -- 69
        46581 => X"46",  -- 70
        46582 => X"46",  -- 70
        46583 => X"45",  -- 69
        46584 => X"42",  -- 66
        46585 => X"42",  -- 66
        46586 => X"45",  -- 69
        46587 => X"49",  -- 73
        46588 => X"4A",  -- 74
        46589 => X"47",  -- 71
        46590 => X"46",  -- 70
        46591 => X"48",  -- 72
        46592 => X"3D",  -- 61
        46593 => X"3E",  -- 62
        46594 => X"3C",  -- 60
        46595 => X"3B",  -- 59
        46596 => X"3E",  -- 62
        46597 => X"41",  -- 65
        46598 => X"3E",  -- 62
        46599 => X"38",  -- 56
        46600 => X"37",  -- 55
        46601 => X"40",  -- 64
        46602 => X"43",  -- 67
        46603 => X"3F",  -- 63
        46604 => X"3D",  -- 61
        46605 => X"42",  -- 66
        46606 => X"43",  -- 67
        46607 => X"40",  -- 64
        46608 => X"3F",  -- 63
        46609 => X"3F",  -- 63
        46610 => X"40",  -- 64
        46611 => X"44",  -- 68
        46612 => X"43",  -- 67
        46613 => X"3E",  -- 62
        46614 => X"3C",  -- 60
        46615 => X"3E",  -- 62
        46616 => X"3C",  -- 60
        46617 => X"42",  -- 66
        46618 => X"47",  -- 71
        46619 => X"43",  -- 67
        46620 => X"3F",  -- 63
        46621 => X"40",  -- 64
        46622 => X"43",  -- 67
        46623 => X"45",  -- 69
        46624 => X"44",  -- 68
        46625 => X"4B",  -- 75
        46626 => X"45",  -- 69
        46627 => X"41",  -- 65
        46628 => X"50",  -- 80
        46629 => X"68",  -- 104
        46630 => X"79",  -- 121
        46631 => X"85",  -- 133
        46632 => X"86",  -- 134
        46633 => X"8A",  -- 138
        46634 => X"93",  -- 147
        46635 => X"92",  -- 146
        46636 => X"9D",  -- 157
        46637 => X"A4",  -- 164
        46638 => X"9E",  -- 158
        46639 => X"AA",  -- 170
        46640 => X"98",  -- 152
        46641 => X"8D",  -- 141
        46642 => X"81",  -- 129
        46643 => X"84",  -- 132
        46644 => X"92",  -- 146
        46645 => X"96",  -- 150
        46646 => X"99",  -- 153
        46647 => X"A5",  -- 165
        46648 => X"A1",  -- 161
        46649 => X"A9",  -- 169
        46650 => X"A0",  -- 160
        46651 => X"AC",  -- 172
        46652 => X"AA",  -- 170
        46653 => X"92",  -- 146
        46654 => X"96",  -- 150
        46655 => X"98",  -- 152
        46656 => X"A0",  -- 160
        46657 => X"98",  -- 152
        46658 => X"A6",  -- 166
        46659 => X"A6",  -- 166
        46660 => X"96",  -- 150
        46661 => X"9A",  -- 154
        46662 => X"A6",  -- 166
        46663 => X"B3",  -- 179
        46664 => X"B6",  -- 182
        46665 => X"B3",  -- 179
        46666 => X"B0",  -- 176
        46667 => X"B3",  -- 179
        46668 => X"B5",  -- 181
        46669 => X"B2",  -- 178
        46670 => X"AF",  -- 175
        46671 => X"A9",  -- 169
        46672 => X"A5",  -- 165
        46673 => X"AC",  -- 172
        46674 => X"AC",  -- 172
        46675 => X"A7",  -- 167
        46676 => X"AA",  -- 170
        46677 => X"B4",  -- 180
        46678 => X"B4",  -- 180
        46679 => X"AC",  -- 172
        46680 => X"B0",  -- 176
        46681 => X"B2",  -- 178
        46682 => X"B6",  -- 182
        46683 => X"BA",  -- 186
        46684 => X"BD",  -- 189
        46685 => X"BE",  -- 190
        46686 => X"BF",  -- 191
        46687 => X"C1",  -- 193
        46688 => X"C9",  -- 201
        46689 => X"CB",  -- 203
        46690 => X"CC",  -- 204
        46691 => X"CB",  -- 203
        46692 => X"C7",  -- 199
        46693 => X"C1",  -- 193
        46694 => X"BB",  -- 187
        46695 => X"B7",  -- 183
        46696 => X"B8",  -- 184
        46697 => X"BD",  -- 189
        46698 => X"BD",  -- 189
        46699 => X"B5",  -- 181
        46700 => X"AE",  -- 174
        46701 => X"A3",  -- 163
        46702 => X"8B",  -- 139
        46703 => X"73",  -- 115
        46704 => X"45",  -- 69
        46705 => X"4F",  -- 79
        46706 => X"72",  -- 114
        46707 => X"5B",  -- 91
        46708 => X"49",  -- 73
        46709 => X"4F",  -- 79
        46710 => X"31",  -- 49
        46711 => X"37",  -- 55
        46712 => X"3E",  -- 62
        46713 => X"4C",  -- 76
        46714 => X"58",  -- 88
        46715 => X"63",  -- 99
        46716 => X"6A",  -- 106
        46717 => X"66",  -- 102
        46718 => X"6C",  -- 108
        46719 => X"7E",  -- 126
        46720 => X"68",  -- 104
        46721 => X"6B",  -- 107
        46722 => X"6C",  -- 108
        46723 => X"6B",  -- 107
        46724 => X"6E",  -- 110
        46725 => X"76",  -- 118
        46726 => X"80",  -- 128
        46727 => X"85",  -- 133
        46728 => X"7F",  -- 127
        46729 => X"83",  -- 131
        46730 => X"89",  -- 137
        46731 => X"8B",  -- 139
        46732 => X"86",  -- 134
        46733 => X"7F",  -- 127
        46734 => X"7C",  -- 124
        46735 => X"7F",  -- 127
        46736 => X"80",  -- 128
        46737 => X"79",  -- 121
        46738 => X"6E",  -- 110
        46739 => X"66",  -- 102
        46740 => X"60",  -- 96
        46741 => X"5A",  -- 90
        46742 => X"55",  -- 85
        46743 => X"51",  -- 81
        46744 => X"55",  -- 85
        46745 => X"55",  -- 85
        46746 => X"57",  -- 87
        46747 => X"54",  -- 84
        46748 => X"53",  -- 83
        46749 => X"54",  -- 84
        46750 => X"58",  -- 88
        46751 => X"5B",  -- 91
        46752 => X"64",  -- 100
        46753 => X"62",  -- 98
        46754 => X"6C",  -- 108
        46755 => X"7B",  -- 123
        46756 => X"7B",  -- 123
        46757 => X"69",  -- 105
        46758 => X"60",  -- 96
        46759 => X"64",  -- 100
        46760 => X"5F",  -- 95
        46761 => X"59",  -- 89
        46762 => X"57",  -- 87
        46763 => X"64",  -- 100
        46764 => X"6B",  -- 107
        46765 => X"55",  -- 85
        46766 => X"29",  -- 41
        46767 => X"04",  -- 4
        46768 => X"01",  -- 1
        46769 => X"0E",  -- 14
        46770 => X"28",  -- 40
        46771 => X"3C",  -- 60
        46772 => X"4C",  -- 76
        46773 => X"5E",  -- 94
        46774 => X"61",  -- 97
        46775 => X"53",  -- 83
        46776 => X"28",  -- 40
        46777 => X"7A",  -- 122
        46778 => X"7B",  -- 123
        46779 => X"3B",  -- 59
        46780 => X"69",  -- 105
        46781 => X"6C",  -- 108
        46782 => X"6E",  -- 110
        46783 => X"50",  -- 80
        46784 => X"43",  -- 67
        46785 => X"68",  -- 104
        46786 => X"5F",  -- 95
        46787 => X"45",  -- 69
        46788 => X"47",  -- 71
        46789 => X"44",  -- 68
        46790 => X"39",  -- 57
        46791 => X"45",  -- 69
        46792 => X"38",  -- 56
        46793 => X"3B",  -- 59
        46794 => X"3B",  -- 59
        46795 => X"38",  -- 56
        46796 => X"3B",  -- 59
        46797 => X"46",  -- 70
        46798 => X"54",  -- 84
        46799 => X"5D",  -- 93
        46800 => X"56",  -- 86
        46801 => X"5F",  -- 95
        46802 => X"5E",  -- 94
        46803 => X"54",  -- 84
        46804 => X"4F",  -- 79
        46805 => X"51",  -- 81
        46806 => X"56",  -- 86
        46807 => X"5B",  -- 91
        46808 => X"5E",  -- 94
        46809 => X"6A",  -- 106
        46810 => X"75",  -- 117
        46811 => X"7C",  -- 124
        46812 => X"83",  -- 131
        46813 => X"87",  -- 135
        46814 => X"80",  -- 128
        46815 => X"74",  -- 116
        46816 => X"7C",  -- 124
        46817 => X"7D",  -- 125
        46818 => X"72",  -- 114
        46819 => X"67",  -- 103
        46820 => X"6D",  -- 109
        46821 => X"73",  -- 115
        46822 => X"77",  -- 119
        46823 => X"7F",  -- 127
        46824 => X"74",  -- 116
        46825 => X"7E",  -- 126
        46826 => X"88",  -- 136
        46827 => X"86",  -- 134
        46828 => X"7E",  -- 126
        46829 => X"77",  -- 119
        46830 => X"71",  -- 113
        46831 => X"6F",  -- 111
        46832 => X"5E",  -- 94
        46833 => X"61",  -- 97
        46834 => X"5C",  -- 92
        46835 => X"56",  -- 86
        46836 => X"5D",  -- 93
        46837 => X"60",  -- 96
        46838 => X"63",  -- 99
        46839 => X"6C",  -- 108
        46840 => X"68",  -- 104
        46841 => X"6D",  -- 109
        46842 => X"7B",  -- 123
        46843 => X"76",  -- 118
        46844 => X"56",  -- 86
        46845 => X"36",  -- 54
        46846 => X"43",  -- 67
        46847 => X"7A",  -- 122
        46848 => X"7A",  -- 122
        46849 => X"71",  -- 113
        46850 => X"BA",  -- 186
        46851 => X"88",  -- 136
        46852 => X"63",  -- 99
        46853 => X"3E",  -- 62
        46854 => X"26",  -- 38
        46855 => X"62",  -- 98
        46856 => X"98",  -- 152
        46857 => X"A7",  -- 167
        46858 => X"91",  -- 145
        46859 => X"6F",  -- 111
        46860 => X"36",  -- 54
        46861 => X"09",  -- 9
        46862 => X"16",  -- 22
        46863 => X"1F",  -- 31
        46864 => X"18",  -- 24
        46865 => X"19",  -- 25
        46866 => X"45",  -- 69
        46867 => X"4D",  -- 77
        46868 => X"46",  -- 70
        46869 => X"37",  -- 55
        46870 => X"23",  -- 35
        46871 => X"4C",  -- 76
        46872 => X"5D",  -- 93
        46873 => X"74",  -- 116
        46874 => X"73",  -- 115
        46875 => X"72",  -- 114
        46876 => X"7F",  -- 127
        46877 => X"78",  -- 120
        46878 => X"84",  -- 132
        46879 => X"8F",  -- 143
        46880 => X"A3",  -- 163
        46881 => X"AA",  -- 170
        46882 => X"AC",  -- 172
        46883 => X"B2",  -- 178
        46884 => X"AD",  -- 173
        46885 => X"B0",  -- 176
        46886 => X"C4",  -- 196
        46887 => X"C1",  -- 193
        46888 => X"C5",  -- 197
        46889 => X"BB",  -- 187
        46890 => X"AC",  -- 172
        46891 => X"A7",  -- 167
        46892 => X"8D",  -- 141
        46893 => X"63",  -- 99
        46894 => X"46",  -- 70
        46895 => X"4D",  -- 77
        46896 => X"49",  -- 73
        46897 => X"47",  -- 71
        46898 => X"44",  -- 68
        46899 => X"42",  -- 66
        46900 => X"41",  -- 65
        46901 => X"43",  -- 67
        46902 => X"45",  -- 69
        46903 => X"46",  -- 70
        46904 => X"44",  -- 68
        46905 => X"42",  -- 66
        46906 => X"45",  -- 69
        46907 => X"49",  -- 73
        46908 => X"49",  -- 73
        46909 => X"45",  -- 69
        46910 => X"42",  -- 66
        46911 => X"43",  -- 67
        46912 => X"3E",  -- 62
        46913 => X"3D",  -- 61
        46914 => X"3B",  -- 59
        46915 => X"3A",  -- 58
        46916 => X"3C",  -- 60
        46917 => X"3E",  -- 62
        46918 => X"3D",  -- 61
        46919 => X"39",  -- 57
        46920 => X"34",  -- 52
        46921 => X"3C",  -- 60
        46922 => X"40",  -- 64
        46923 => X"3D",  -- 61
        46924 => X"3B",  -- 59
        46925 => X"3F",  -- 63
        46926 => X"40",  -- 64
        46927 => X"3D",  -- 61
        46928 => X"3D",  -- 61
        46929 => X"3D",  -- 61
        46930 => X"3F",  -- 63
        46931 => X"43",  -- 67
        46932 => X"44",  -- 68
        46933 => X"40",  -- 64
        46934 => X"3D",  -- 61
        46935 => X"3D",  -- 61
        46936 => X"3D",  -- 61
        46937 => X"3F",  -- 63
        46938 => X"44",  -- 68
        46939 => X"46",  -- 70
        46940 => X"42",  -- 66
        46941 => X"3E",  -- 62
        46942 => X"40",  -- 64
        46943 => X"44",  -- 68
        46944 => X"46",  -- 70
        46945 => X"4B",  -- 75
        46946 => X"47",  -- 71
        46947 => X"48",  -- 72
        46948 => X"5C",  -- 92
        46949 => X"70",  -- 112
        46950 => X"7D",  -- 125
        46951 => X"86",  -- 134
        46952 => X"7E",  -- 126
        46953 => X"81",  -- 129
        46954 => X"8D",  -- 141
        46955 => X"8E",  -- 142
        46956 => X"9C",  -- 156
        46957 => X"A6",  -- 166
        46958 => X"A1",  -- 161
        46959 => X"AD",  -- 173
        46960 => X"9C",  -- 156
        46961 => X"9B",  -- 155
        46962 => X"85",  -- 133
        46963 => X"71",  -- 113
        46964 => X"82",  -- 130
        46965 => X"9F",  -- 159
        46966 => X"A8",  -- 168
        46967 => X"A3",  -- 163
        46968 => X"98",  -- 152
        46969 => X"A4",  -- 164
        46970 => X"9A",  -- 154
        46971 => X"AF",  -- 175
        46972 => X"AC",  -- 172
        46973 => X"94",  -- 148
        46974 => X"A4",  -- 164
        46975 => X"A1",  -- 161
        46976 => X"A6",  -- 166
        46977 => X"A3",  -- 163
        46978 => X"A2",  -- 162
        46979 => X"AB",  -- 171
        46980 => X"A0",  -- 160
        46981 => X"99",  -- 153
        46982 => X"A5",  -- 165
        46983 => X"A5",  -- 165
        46984 => X"AD",  -- 173
        46985 => X"B5",  -- 181
        46986 => X"A9",  -- 169
        46987 => X"B2",  -- 178
        46988 => X"B5",  -- 181
        46989 => X"AE",  -- 174
        46990 => X"B7",  -- 183
        46991 => X"AC",  -- 172
        46992 => X"A5",  -- 165
        46993 => X"AC",  -- 172
        46994 => X"AF",  -- 175
        46995 => X"AE",  -- 174
        46996 => X"AF",  -- 175
        46997 => X"B2",  -- 178
        46998 => X"B4",  -- 180
        46999 => X"B5",  -- 181
        47000 => X"B5",  -- 181
        47001 => X"B5",  -- 181
        47002 => X"B7",  -- 183
        47003 => X"B9",  -- 185
        47004 => X"BE",  -- 190
        47005 => X"C1",  -- 193
        47006 => X"C1",  -- 193
        47007 => X"C1",  -- 193
        47008 => X"C7",  -- 199
        47009 => X"CA",  -- 202
        47010 => X"CE",  -- 206
        47011 => X"CD",  -- 205
        47012 => X"C8",  -- 200
        47013 => X"C2",  -- 194
        47014 => X"BD",  -- 189
        47015 => X"BC",  -- 188
        47016 => X"B3",  -- 179
        47017 => X"B9",  -- 185
        47018 => X"BD",  -- 189
        47019 => X"B8",  -- 184
        47020 => X"B0",  -- 176
        47021 => X"A5",  -- 165
        47022 => X"94",  -- 148
        47023 => X"86",  -- 134
        47024 => X"63",  -- 99
        47025 => X"4E",  -- 78
        47026 => X"3F",  -- 63
        47027 => X"4E",  -- 78
        47028 => X"4B",  -- 75
        47029 => X"38",  -- 56
        47030 => X"3A",  -- 58
        47031 => X"48",  -- 72
        47032 => X"3F",  -- 63
        47033 => X"45",  -- 69
        47034 => X"4D",  -- 77
        47035 => X"5C",  -- 92
        47036 => X"6A",  -- 106
        47037 => X"6B",  -- 107
        47038 => X"6E",  -- 110
        47039 => X"7A",  -- 122
        47040 => X"70",  -- 112
        47041 => X"74",  -- 116
        47042 => X"76",  -- 118
        47043 => X"76",  -- 118
        47044 => X"75",  -- 117
        47045 => X"76",  -- 118
        47046 => X"7B",  -- 123
        47047 => X"7E",  -- 126
        47048 => X"79",  -- 121
        47049 => X"7E",  -- 126
        47050 => X"83",  -- 131
        47051 => X"83",  -- 131
        47052 => X"7E",  -- 126
        47053 => X"79",  -- 121
        47054 => X"7A",  -- 122
        47055 => X"7D",  -- 125
        47056 => X"81",  -- 129
        47057 => X"7A",  -- 122
        47058 => X"70",  -- 112
        47059 => X"67",  -- 103
        47060 => X"60",  -- 96
        47061 => X"5C",  -- 92
        47062 => X"57",  -- 87
        47063 => X"53",  -- 83
        47064 => X"4F",  -- 79
        47065 => X"4E",  -- 78
        47066 => X"4D",  -- 77
        47067 => X"4C",  -- 76
        47068 => X"4A",  -- 74
        47069 => X"4B",  -- 75
        47070 => X"4D",  -- 77
        47071 => X"50",  -- 80
        47072 => X"5F",  -- 95
        47073 => X"5C",  -- 92
        47074 => X"6D",  -- 109
        47075 => X"80",  -- 128
        47076 => X"76",  -- 118
        47077 => X"63",  -- 99
        47078 => X"5F",  -- 95
        47079 => X"68",  -- 104
        47080 => X"5C",  -- 92
        47081 => X"61",  -- 97
        47082 => X"63",  -- 99
        47083 => X"6A",  -- 106
        47084 => X"61",  -- 97
        47085 => X"4D",  -- 77
        47086 => X"38",  -- 56
        47087 => X"1C",  -- 28
        47088 => X"06",  -- 6
        47089 => X"09",  -- 9
        47090 => X"12",  -- 18
        47091 => X"1C",  -- 28
        47092 => X"2D",  -- 45
        47093 => X"49",  -- 73
        47094 => X"5D",  -- 93
        47095 => X"5A",  -- 90
        47096 => X"53",  -- 83
        47097 => X"77",  -- 119
        47098 => X"72",  -- 114
        47099 => X"51",  -- 81
        47100 => X"77",  -- 119
        47101 => X"6C",  -- 108
        47102 => X"50",  -- 80
        47103 => X"1B",  -- 27
        47104 => X"41",  -- 65
        47105 => X"66",  -- 102
        47106 => X"5B",  -- 91
        47107 => X"39",  -- 57
        47108 => X"3B",  -- 59
        47109 => X"3F",  -- 63
        47110 => X"37",  -- 55
        47111 => X"3E",  -- 62
        47112 => X"33",  -- 51
        47113 => X"31",  -- 49
        47114 => X"2E",  -- 46
        47115 => X"2F",  -- 47
        47116 => X"37",  -- 55
        47117 => X"41",  -- 65
        47118 => X"4A",  -- 74
        47119 => X"50",  -- 80
        47120 => X"5E",  -- 94
        47121 => X"52",  -- 82
        47122 => X"58",  -- 88
        47123 => X"5D",  -- 93
        47124 => X"5A",  -- 90
        47125 => X"68",  -- 104
        47126 => X"6F",  -- 111
        47127 => X"5C",  -- 92
        47128 => X"61",  -- 97
        47129 => X"69",  -- 105
        47130 => X"71",  -- 113
        47131 => X"77",  -- 119
        47132 => X"82",  -- 130
        47133 => X"8B",  -- 139
        47134 => X"88",  -- 136
        47135 => X"7E",  -- 126
        47136 => X"7B",  -- 123
        47137 => X"82",  -- 130
        47138 => X"7E",  -- 126
        47139 => X"79",  -- 121
        47140 => X"7F",  -- 127
        47141 => X"7F",  -- 127
        47142 => X"7B",  -- 123
        47143 => X"7E",  -- 126
        47144 => X"7A",  -- 122
        47145 => X"7E",  -- 126
        47146 => X"82",  -- 130
        47147 => X"7F",  -- 127
        47148 => X"76",  -- 118
        47149 => X"6E",  -- 110
        47150 => X"67",  -- 103
        47151 => X"64",  -- 100
        47152 => X"67",  -- 103
        47153 => X"5A",  -- 90
        47154 => X"4B",  -- 75
        47155 => X"4E",  -- 78
        47156 => X"62",  -- 98
        47157 => X"6A",  -- 106
        47158 => X"6C",  -- 108
        47159 => X"70",  -- 112
        47160 => X"6B",  -- 107
        47161 => X"5C",  -- 92
        47162 => X"72",  -- 114
        47163 => X"82",  -- 130
        47164 => X"78",  -- 120
        47165 => X"50",  -- 80
        47166 => X"3A",  -- 58
        47167 => X"6C",  -- 108
        47168 => X"8B",  -- 139
        47169 => X"85",  -- 133
        47170 => X"BA",  -- 186
        47171 => X"C7",  -- 199
        47172 => X"A0",  -- 160
        47173 => X"68",  -- 104
        47174 => X"7D",  -- 125
        47175 => X"A5",  -- 165
        47176 => X"9E",  -- 158
        47177 => X"9F",  -- 159
        47178 => X"7D",  -- 125
        47179 => X"52",  -- 82
        47180 => X"2F",  -- 47
        47181 => X"1D",  -- 29
        47182 => X"23",  -- 35
        47183 => X"1A",  -- 26
        47184 => X"1A",  -- 26
        47185 => X"2F",  -- 47
        47186 => X"56",  -- 86
        47187 => X"3D",  -- 61
        47188 => X"28",  -- 40
        47189 => X"2D",  -- 45
        47190 => X"26",  -- 38
        47191 => X"4C",  -- 76
        47192 => X"6A",  -- 106
        47193 => X"77",  -- 119
        47194 => X"7A",  -- 122
        47195 => X"74",  -- 116
        47196 => X"7E",  -- 126
        47197 => X"71",  -- 113
        47198 => X"8A",  -- 138
        47199 => X"94",  -- 148
        47200 => X"A1",  -- 161
        47201 => X"A8",  -- 168
        47202 => X"AB",  -- 171
        47203 => X"B3",  -- 179
        47204 => X"AE",  -- 174
        47205 => X"AF",  -- 175
        47206 => X"C2",  -- 194
        47207 => X"BF",  -- 191
        47208 => X"C6",  -- 198
        47209 => X"C1",  -- 193
        47210 => X"A8",  -- 168
        47211 => X"9A",  -- 154
        47212 => X"7B",  -- 123
        47213 => X"72",  -- 114
        47214 => X"53",  -- 83
        47215 => X"3F",  -- 63
        47216 => X"47",  -- 71
        47217 => X"45",  -- 69
        47218 => X"42",  -- 66
        47219 => X"3F",  -- 63
        47220 => X"3E",  -- 62
        47221 => X"3F",  -- 63
        47222 => X"42",  -- 66
        47223 => X"45",  -- 69
        47224 => X"44",  -- 68
        47225 => X"43",  -- 67
        47226 => X"45",  -- 69
        47227 => X"49",  -- 73
        47228 => X"49",  -- 73
        47229 => X"44",  -- 68
        47230 => X"40",  -- 64
        47231 => X"3F",  -- 63
        47232 => X"3E",  -- 62
        47233 => X"3C",  -- 60
        47234 => X"3A",  -- 58
        47235 => X"38",  -- 56
        47236 => X"39",  -- 57
        47237 => X"3B",  -- 59
        47238 => X"3B",  -- 59
        47239 => X"3A",  -- 58
        47240 => X"32",  -- 50
        47241 => X"39",  -- 57
        47242 => X"3D",  -- 61
        47243 => X"3B",  -- 59
        47244 => X"3A",  -- 58
        47245 => X"3C",  -- 60
        47246 => X"3D",  -- 61
        47247 => X"3B",  -- 59
        47248 => X"3D",  -- 61
        47249 => X"3C",  -- 60
        47250 => X"3F",  -- 63
        47251 => X"42",  -- 66
        47252 => X"43",  -- 67
        47253 => X"42",  -- 66
        47254 => X"3F",  -- 63
        47255 => X"3D",  -- 61
        47256 => X"3E",  -- 62
        47257 => X"3D",  -- 61
        47258 => X"42",  -- 66
        47259 => X"47",  -- 71
        47260 => X"45",  -- 69
        47261 => X"3D",  -- 61
        47262 => X"3E",  -- 62
        47263 => X"45",  -- 69
        47264 => X"49",  -- 73
        47265 => X"4B",  -- 75
        47266 => X"49",  -- 73
        47267 => X"50",  -- 80
        47268 => X"66",  -- 102
        47269 => X"77",  -- 119
        47270 => X"7D",  -- 125
        47271 => X"82",  -- 130
        47272 => X"7D",  -- 125
        47273 => X"7F",  -- 127
        47274 => X"8A",  -- 138
        47275 => X"8C",  -- 140
        47276 => X"9A",  -- 154
        47277 => X"A6",  -- 166
        47278 => X"A1",  -- 161
        47279 => X"AC",  -- 172
        47280 => X"A6",  -- 166
        47281 => X"A2",  -- 162
        47282 => X"82",  -- 130
        47283 => X"66",  -- 102
        47284 => X"7A",  -- 122
        47285 => X"A3",  -- 163
        47286 => X"AB",  -- 171
        47287 => X"9D",  -- 157
        47288 => X"95",  -- 149
        47289 => X"A2",  -- 162
        47290 => X"97",  -- 151
        47291 => X"AE",  -- 174
        47292 => X"A9",  -- 169
        47293 => X"96",  -- 150
        47294 => X"B2",  -- 178
        47295 => X"AD",  -- 173
        47296 => X"AD",  -- 173
        47297 => X"AC",  -- 172
        47298 => X"9F",  -- 159
        47299 => X"AB",  -- 171
        47300 => X"A8",  -- 168
        47301 => X"9A",  -- 154
        47302 => X"A5",  -- 165
        47303 => X"9F",  -- 159
        47304 => X"A4",  -- 164
        47305 => X"B5",  -- 181
        47306 => X"A4",  -- 164
        47307 => X"B1",  -- 177
        47308 => X"B5",  -- 181
        47309 => X"AC",  -- 172
        47310 => X"C0",  -- 192
        47311 => X"B0",  -- 176
        47312 => X"B0",  -- 176
        47313 => X"B0",  -- 176
        47314 => X"B2",  -- 178
        47315 => X"B6",  -- 182
        47316 => X"B6",  -- 182
        47317 => X"B5",  -- 181
        47318 => X"B6",  -- 182
        47319 => X"B9",  -- 185
        47320 => X"BC",  -- 188
        47321 => X"BA",  -- 186
        47322 => X"B7",  -- 183
        47323 => X"BA",  -- 186
        47324 => X"BF",  -- 191
        47325 => X"C1",  -- 193
        47326 => X"C3",  -- 195
        47327 => X"C2",  -- 194
        47328 => X"C4",  -- 196
        47329 => X"C9",  -- 201
        47330 => X"CE",  -- 206
        47331 => X"CE",  -- 206
        47332 => X"C8",  -- 200
        47333 => X"C3",  -- 195
        47334 => X"C0",  -- 192
        47335 => X"C0",  -- 192
        47336 => X"B2",  -- 178
        47337 => X"B3",  -- 179
        47338 => X"B3",  -- 179
        47339 => X"B3",  -- 179
        47340 => X"B0",  -- 176
        47341 => X"A7",  -- 167
        47342 => X"97",  -- 151
        47343 => X"8A",  -- 138
        47344 => X"79",  -- 121
        47345 => X"59",  -- 89
        47346 => X"32",  -- 50
        47347 => X"50",  -- 80
        47348 => X"54",  -- 84
        47349 => X"2F",  -- 47
        47350 => X"36",  -- 54
        47351 => X"39",  -- 57
        47352 => X"44",  -- 68
        47353 => X"45",  -- 69
        47354 => X"48",  -- 72
        47355 => X"55",  -- 85
        47356 => X"66",  -- 102
        47357 => X"6A",  -- 106
        47358 => X"70",  -- 112
        47359 => X"7C",  -- 124
        47360 => X"73",  -- 115
        47361 => X"78",  -- 120
        47362 => X"80",  -- 128
        47363 => X"84",  -- 132
        47364 => X"83",  -- 131
        47365 => X"7F",  -- 127
        47366 => X"7B",  -- 123
        47367 => X"7B",  -- 123
        47368 => X"77",  -- 119
        47369 => X"7C",  -- 124
        47370 => X"7D",  -- 125
        47371 => X"79",  -- 121
        47372 => X"74",  -- 116
        47373 => X"73",  -- 115
        47374 => X"77",  -- 119
        47375 => X"7B",  -- 123
        47376 => X"7C",  -- 124
        47377 => X"79",  -- 121
        47378 => X"72",  -- 114
        47379 => X"6B",  -- 107
        47380 => X"62",  -- 98
        47381 => X"5D",  -- 93
        47382 => X"57",  -- 87
        47383 => X"54",  -- 84
        47384 => X"4D",  -- 77
        47385 => X"4B",  -- 75
        47386 => X"48",  -- 72
        47387 => X"45",  -- 69
        47388 => X"45",  -- 69
        47389 => X"46",  -- 70
        47390 => X"49",  -- 73
        47391 => X"4B",  -- 75
        47392 => X"54",  -- 84
        47393 => X"56",  -- 86
        47394 => X"70",  -- 112
        47395 => X"82",  -- 130
        47396 => X"70",  -- 112
        47397 => X"5B",  -- 91
        47398 => X"5F",  -- 95
        47399 => X"69",  -- 105
        47400 => X"5A",  -- 90
        47401 => X"64",  -- 100
        47402 => X"67",  -- 103
        47403 => X"6B",  -- 107
        47404 => X"5B",  -- 91
        47405 => X"4C",  -- 76
        47406 => X"4B",  -- 75
        47407 => X"32",  -- 50
        47408 => X"0D",  -- 13
        47409 => X"08",  -- 8
        47410 => X"08",  -- 8
        47411 => X"0E",  -- 14
        47412 => X"1F",  -- 31
        47413 => X"3B",  -- 59
        47414 => X"4F",  -- 79
        47415 => X"4C",  -- 76
        47416 => X"5C",  -- 92
        47417 => X"6F",  -- 111
        47418 => X"59",  -- 89
        47419 => X"3F",  -- 63
        47420 => X"6C",  -- 108
        47421 => X"79",  -- 121
        47422 => X"45",  -- 69
        47423 => X"28",  -- 40
        47424 => X"5B",  -- 91
        47425 => X"63",  -- 99
        47426 => X"59",  -- 89
        47427 => X"43",  -- 67
        47428 => X"3A",  -- 58
        47429 => X"3D",  -- 61
        47430 => X"40",  -- 64
        47431 => X"39",  -- 57
        47432 => X"37",  -- 55
        47433 => X"31",  -- 49
        47434 => X"2C",  -- 44
        47435 => X"30",  -- 48
        47436 => X"39",  -- 57
        47437 => X"42",  -- 66
        47438 => X"48",  -- 72
        47439 => X"4A",  -- 74
        47440 => X"43",  -- 67
        47441 => X"4C",  -- 76
        47442 => X"44",  -- 68
        47443 => X"4B",  -- 75
        47444 => X"69",  -- 105
        47445 => X"6E",  -- 110
        47446 => X"61",  -- 97
        47447 => X"62",  -- 98
        47448 => X"70",  -- 112
        47449 => X"72",  -- 114
        47450 => X"72",  -- 114
        47451 => X"72",  -- 114
        47452 => X"7C",  -- 124
        47453 => X"88",  -- 136
        47454 => X"8C",  -- 140
        47455 => X"87",  -- 135
        47456 => X"77",  -- 119
        47457 => X"7F",  -- 127
        47458 => X"7D",  -- 125
        47459 => X"7A",  -- 122
        47460 => X"7D",  -- 125
        47461 => X"7E",  -- 126
        47462 => X"78",  -- 120
        47463 => X"79",  -- 121
        47464 => X"80",  -- 128
        47465 => X"7A",  -- 122
        47466 => X"75",  -- 117
        47467 => X"70",  -- 112
        47468 => X"6C",  -- 108
        47469 => X"69",  -- 105
        47470 => X"68",  -- 104
        47471 => X"67",  -- 103
        47472 => X"67",  -- 103
        47473 => X"5B",  -- 91
        47474 => X"4A",  -- 74
        47475 => X"4D",  -- 77
        47476 => X"62",  -- 98
        47477 => X"6E",  -- 110
        47478 => X"70",  -- 112
        47479 => X"76",  -- 118
        47480 => X"6D",  -- 109
        47481 => X"64",  -- 100
        47482 => X"6E",  -- 110
        47483 => X"7A",  -- 122
        47484 => X"8E",  -- 142
        47485 => X"84",  -- 132
        47486 => X"67",  -- 103
        47487 => X"7F",  -- 127
        47488 => X"9C",  -- 156
        47489 => X"A1",  -- 161
        47490 => X"CB",  -- 203
        47491 => X"E3",  -- 227
        47492 => X"D6",  -- 214
        47493 => X"C4",  -- 196
        47494 => X"D0",  -- 208
        47495 => X"B7",  -- 183
        47496 => X"A8",  -- 168
        47497 => X"89",  -- 137
        47498 => X"58",  -- 88
        47499 => X"41",  -- 65
        47500 => X"42",  -- 66
        47501 => X"48",  -- 72
        47502 => X"46",  -- 70
        47503 => X"34",  -- 52
        47504 => X"18",  -- 24
        47505 => X"33",  -- 51
        47506 => X"40",  -- 64
        47507 => X"2C",  -- 44
        47508 => X"1D",  -- 29
        47509 => X"22",  -- 34
        47510 => X"36",  -- 54
        47511 => X"53",  -- 83
        47512 => X"75",  -- 117
        47513 => X"7E",  -- 126
        47514 => X"7E",  -- 126
        47515 => X"77",  -- 119
        47516 => X"80",  -- 128
        47517 => X"70",  -- 112
        47518 => X"8A",  -- 138
        47519 => X"99",  -- 153
        47520 => X"A0",  -- 160
        47521 => X"A7",  -- 167
        47522 => X"AB",  -- 171
        47523 => X"B4",  -- 180
        47524 => X"AE",  -- 174
        47525 => X"AC",  -- 172
        47526 => X"BF",  -- 191
        47527 => X"C0",  -- 192
        47528 => X"C2",  -- 194
        47529 => X"B7",  -- 183
        47530 => X"AD",  -- 173
        47531 => X"9E",  -- 158
        47532 => X"68",  -- 104
        47533 => X"67",  -- 103
        47534 => X"59",  -- 89
        47535 => X"3A",  -- 58
        47536 => X"43",  -- 67
        47537 => X"42",  -- 66
        47538 => X"41",  -- 65
        47539 => X"3E",  -- 62
        47540 => X"3B",  -- 59
        47541 => X"3C",  -- 60
        47542 => X"40",  -- 64
        47543 => X"42",  -- 66
        47544 => X"40",  -- 64
        47545 => X"3F",  -- 63
        47546 => X"42",  -- 66
        47547 => X"49",  -- 73
        47548 => X"4A",  -- 74
        47549 => X"46",  -- 70
        47550 => X"40",  -- 64
        47551 => X"3E",  -- 62
        47552 => X"3E",  -- 62
        47553 => X"3B",  -- 59
        47554 => X"38",  -- 56
        47555 => X"37",  -- 55
        47556 => X"37",  -- 55
        47557 => X"38",  -- 56
        47558 => X"39",  -- 57
        47559 => X"3A",  -- 58
        47560 => X"32",  -- 50
        47561 => X"38",  -- 56
        47562 => X"3B",  -- 59
        47563 => X"3B",  -- 59
        47564 => X"39",  -- 57
        47565 => X"3A",  -- 58
        47566 => X"3B",  -- 59
        47567 => X"3B",  -- 59
        47568 => X"3B",  -- 59
        47569 => X"3B",  -- 59
        47570 => X"3C",  -- 60
        47571 => X"3E",  -- 62
        47572 => X"42",  -- 66
        47573 => X"43",  -- 67
        47574 => X"42",  -- 66
        47575 => X"3F",  -- 63
        47576 => X"40",  -- 64
        47577 => X"3E",  -- 62
        47578 => X"40",  -- 64
        47579 => X"46",  -- 70
        47580 => X"45",  -- 69
        47581 => X"3F",  -- 63
        47582 => X"3F",  -- 63
        47583 => X"44",  -- 68
        47584 => X"45",  -- 69
        47585 => X"48",  -- 72
        47586 => X"48",  -- 72
        47587 => X"57",  -- 87
        47588 => X"70",  -- 112
        47589 => X"7D",  -- 125
        47590 => X"7E",  -- 126
        47591 => X"82",  -- 130
        47592 => X"8A",  -- 138
        47593 => X"8A",  -- 138
        47594 => X"8F",  -- 143
        47595 => X"8F",  -- 143
        47596 => X"9C",  -- 156
        47597 => X"A3",  -- 163
        47598 => X"9C",  -- 156
        47599 => X"A7",  -- 167
        47600 => X"A7",  -- 167
        47601 => X"A5",  -- 165
        47602 => X"8B",  -- 139
        47603 => X"70",  -- 112
        47604 => X"7A",  -- 122
        47605 => X"93",  -- 147
        47606 => X"9F",  -- 159
        47607 => X"9F",  -- 159
        47608 => X"A1",  -- 161
        47609 => X"A7",  -- 167
        47610 => X"9F",  -- 159
        47611 => X"AF",  -- 175
        47612 => X"A6",  -- 166
        47613 => X"9A",  -- 154
        47614 => X"B8",  -- 184
        47615 => X"B4",  -- 180
        47616 => X"B1",  -- 177
        47617 => X"B1",  -- 177
        47618 => X"9E",  -- 158
        47619 => X"A7",  -- 167
        47620 => X"AA",  -- 170
        47621 => X"9C",  -- 156
        47622 => X"A5",  -- 165
        47623 => X"A2",  -- 162
        47624 => X"9E",  -- 158
        47625 => X"B1",  -- 177
        47626 => X"A2",  -- 162
        47627 => X"B0",  -- 176
        47628 => X"B3",  -- 179
        47629 => X"AE",  -- 174
        47630 => X"C6",  -- 198
        47631 => X"B8",  -- 184
        47632 => X"B6",  -- 182
        47633 => X"B1",  -- 177
        47634 => X"B1",  -- 177
        47635 => X"B6",  -- 182
        47636 => X"BA",  -- 186
        47637 => X"BA",  -- 186
        47638 => X"BB",  -- 187
        47639 => X"BF",  -- 191
        47640 => X"BE",  -- 190
        47641 => X"BB",  -- 187
        47642 => X"BA",  -- 186
        47643 => X"BC",  -- 188
        47644 => X"C0",  -- 192
        47645 => X"C2",  -- 194
        47646 => X"C3",  -- 195
        47647 => X"C2",  -- 194
        47648 => X"C1",  -- 193
        47649 => X"C8",  -- 200
        47650 => X"CE",  -- 206
        47651 => X"CE",  -- 206
        47652 => X"C9",  -- 201
        47653 => X"C4",  -- 196
        47654 => X"C2",  -- 194
        47655 => X"C2",  -- 194
        47656 => X"B5",  -- 181
        47657 => X"AF",  -- 175
        47658 => X"A8",  -- 168
        47659 => X"A9",  -- 169
        47660 => X"B0",  -- 176
        47661 => X"AF",  -- 175
        47662 => X"9D",  -- 157
        47663 => X"89",  -- 137
        47664 => X"7F",  -- 127
        47665 => X"5D",  -- 93
        47666 => X"4F",  -- 79
        47667 => X"30",  -- 48
        47668 => X"32",  -- 50
        47669 => X"47",  -- 71
        47670 => X"32",  -- 50
        47671 => X"33",  -- 51
        47672 => X"3F",  -- 63
        47673 => X"41",  -- 65
        47674 => X"44",  -- 68
        47675 => X"51",  -- 81
        47676 => X"64",  -- 100
        47677 => X"6E",  -- 110
        47678 => X"7A",  -- 122
        47679 => X"8E",  -- 142
        47680 => X"70",  -- 112
        47681 => X"74",  -- 116
        47682 => X"7D",  -- 125
        47683 => X"86",  -- 134
        47684 => X"89",  -- 137
        47685 => X"84",  -- 132
        47686 => X"7E",  -- 126
        47687 => X"7B",  -- 123
        47688 => X"7C",  -- 124
        47689 => X"7E",  -- 126
        47690 => X"7C",  -- 124
        47691 => X"75",  -- 117
        47692 => X"6F",  -- 111
        47693 => X"70",  -- 112
        47694 => X"74",  -- 116
        47695 => X"77",  -- 119
        47696 => X"77",  -- 119
        47697 => X"76",  -- 118
        47698 => X"72",  -- 114
        47699 => X"6E",  -- 110
        47700 => X"65",  -- 101
        47701 => X"5C",  -- 92
        47702 => X"54",  -- 84
        47703 => X"50",  -- 80
        47704 => X"4C",  -- 76
        47705 => X"4A",  -- 74
        47706 => X"47",  -- 71
        47707 => X"45",  -- 69
        47708 => X"44",  -- 68
        47709 => X"44",  -- 68
        47710 => X"47",  -- 71
        47711 => X"47",  -- 71
        47712 => X"4C",  -- 76
        47713 => X"50",  -- 80
        47714 => X"6D",  -- 109
        47715 => X"7E",  -- 126
        47716 => X"67",  -- 103
        47717 => X"55",  -- 85
        47718 => X"5E",  -- 94
        47719 => X"67",  -- 103
        47720 => X"5E",  -- 94
        47721 => X"67",  -- 103
        47722 => X"64",  -- 100
        47723 => X"6C",  -- 108
        47724 => X"5E",  -- 94
        47725 => X"54",  -- 84
        47726 => X"58",  -- 88
        47727 => X"35",  -- 53
        47728 => X"0A",  -- 10
        47729 => X"05",  -- 5
        47730 => X"07",  -- 7
        47731 => X"11",  -- 17
        47732 => X"1F",  -- 31
        47733 => X"34",  -- 52
        47734 => X"40",  -- 64
        47735 => X"39",  -- 57
        47736 => X"4B",  -- 75
        47737 => X"65",  -- 101
        47738 => X"3F",  -- 63
        47739 => X"35",  -- 53
        47740 => X"70",  -- 112
        47741 => X"61",  -- 97
        47742 => X"26",  -- 38
        47743 => X"53",  -- 83
        47744 => X"64",  -- 100
        47745 => X"53",  -- 83
        47746 => X"50",  -- 80
        47747 => X"4B",  -- 75
        47748 => X"3F",  -- 63
        47749 => X"45",  -- 69
        47750 => X"4D",  -- 77
        47751 => X"3E",  -- 62
        47752 => X"43",  -- 67
        47753 => X"3B",  -- 59
        47754 => X"34",  -- 52
        47755 => X"39",  -- 57
        47756 => X"42",  -- 66
        47757 => X"49",  -- 73
        47758 => X"4B",  -- 75
        47759 => X"4C",  -- 76
        47760 => X"4A",  -- 74
        47761 => X"4A",  -- 74
        47762 => X"54",  -- 84
        47763 => X"66",  -- 102
        47764 => X"6F",  -- 111
        47765 => X"70",  -- 112
        47766 => X"71",  -- 113
        47767 => X"70",  -- 112
        47768 => X"7B",  -- 123
        47769 => X"7D",  -- 125
        47770 => X"7A",  -- 122
        47771 => X"77",  -- 119
        47772 => X"7C",  -- 124
        47773 => X"87",  -- 135
        47774 => X"8A",  -- 138
        47775 => X"87",  -- 135
        47776 => X"7F",  -- 127
        47777 => X"82",  -- 130
        47778 => X"7A",  -- 122
        47779 => X"72",  -- 114
        47780 => X"76",  -- 118
        47781 => X"7A",  -- 122
        47782 => X"7B",  -- 123
        47783 => X"80",  -- 128
        47784 => X"7D",  -- 125
        47785 => X"7A",  -- 122
        47786 => X"7D",  -- 125
        47787 => X"82",  -- 130
        47788 => X"80",  -- 128
        47789 => X"76",  -- 118
        47790 => X"69",  -- 105
        47791 => X"60",  -- 96
        47792 => X"62",  -- 98
        47793 => X"64",  -- 100
        47794 => X"5B",  -- 91
        47795 => X"55",  -- 85
        47796 => X"5E",  -- 94
        47797 => X"66",  -- 102
        47798 => X"6E",  -- 110
        47799 => X"7B",  -- 123
        47800 => X"69",  -- 105
        47801 => X"78",  -- 120
        47802 => X"74",  -- 116
        47803 => X"69",  -- 105
        47804 => X"88",  -- 136
        47805 => X"A0",  -- 160
        47806 => X"A0",  -- 160
        47807 => X"AF",  -- 175
        47808 => X"95",  -- 149
        47809 => X"84",  -- 132
        47810 => X"C0",  -- 192
        47811 => X"E0",  -- 224
        47812 => X"E2",  -- 226
        47813 => X"E7",  -- 231
        47814 => X"D2",  -- 210
        47815 => X"BB",  -- 187
        47816 => X"A3",  -- 163
        47817 => X"81",  -- 129
        47818 => X"64",  -- 100
        47819 => X"5A",  -- 90
        47820 => X"4C",  -- 76
        47821 => X"36",  -- 54
        47822 => X"2B",  -- 43
        47823 => X"31",  -- 49
        47824 => X"15",  -- 21
        47825 => X"1F",  -- 31
        47826 => X"19",  -- 25
        47827 => X"23",  -- 35
        47828 => X"26",  -- 38
        47829 => X"21",  -- 33
        47830 => X"42",  -- 66
        47831 => X"5E",  -- 94
        47832 => X"7A",  -- 122
        47833 => X"87",  -- 135
        47834 => X"80",  -- 128
        47835 => X"7E",  -- 126
        47836 => X"85",  -- 133
        47837 => X"73",  -- 115
        47838 => X"80",  -- 128
        47839 => X"96",  -- 150
        47840 => X"A0",  -- 160
        47841 => X"A9",  -- 169
        47842 => X"AF",  -- 175
        47843 => X"B7",  -- 183
        47844 => X"AD",  -- 173
        47845 => X"A8",  -- 168
        47846 => X"BD",  -- 189
        47847 => X"C1",  -- 193
        47848 => X"BC",  -- 188
        47849 => X"A1",  -- 161
        47850 => X"A9",  -- 169
        47851 => X"A8",  -- 168
        47852 => X"64",  -- 100
        47853 => X"46",  -- 70
        47854 => X"48",  -- 72
        47855 => X"40",  -- 64
        47856 => X"3E",  -- 62
        47857 => X"3F",  -- 63
        47858 => X"3E",  -- 62
        47859 => X"3B",  -- 59
        47860 => X"38",  -- 56
        47861 => X"38",  -- 56
        47862 => X"3C",  -- 60
        47863 => X"3F",  -- 63
        47864 => X"3B",  -- 59
        47865 => X"3B",  -- 59
        47866 => X"3F",  -- 63
        47867 => X"47",  -- 71
        47868 => X"4A",  -- 74
        47869 => X"47",  -- 71
        47870 => X"40",  -- 64
        47871 => X"3E",  -- 62
        47872 => X"3D",  -- 61
        47873 => X"3A",  -- 58
        47874 => X"37",  -- 55
        47875 => X"37",  -- 55
        47876 => X"37",  -- 55
        47877 => X"35",  -- 53
        47878 => X"36",  -- 54
        47879 => X"39",  -- 57
        47880 => X"33",  -- 51
        47881 => X"37",  -- 55
        47882 => X"39",  -- 57
        47883 => X"39",  -- 57
        47884 => X"38",  -- 56
        47885 => X"38",  -- 56
        47886 => X"3A",  -- 58
        47887 => X"3C",  -- 60
        47888 => X"3B",  -- 59
        47889 => X"3B",  -- 59
        47890 => X"3A",  -- 58
        47891 => X"3B",  -- 59
        47892 => X"40",  -- 64
        47893 => X"44",  -- 68
        47894 => X"44",  -- 68
        47895 => X"41",  -- 65
        47896 => X"41",  -- 65
        47897 => X"41",  -- 65
        47898 => X"42",  -- 66
        47899 => X"44",  -- 68
        47900 => X"44",  -- 68
        47901 => X"41",  -- 65
        47902 => X"41",  -- 65
        47903 => X"43",  -- 67
        47904 => X"41",  -- 65
        47905 => X"43",  -- 67
        47906 => X"4A",  -- 74
        47907 => X"60",  -- 96
        47908 => X"7C",  -- 124
        47909 => X"84",  -- 132
        47910 => X"83",  -- 131
        47911 => X"88",  -- 136
        47912 => X"92",  -- 146
        47913 => X"90",  -- 144
        47914 => X"91",  -- 145
        47915 => X"8D",  -- 141
        47916 => X"96",  -- 150
        47917 => X"9E",  -- 158
        47918 => X"96",  -- 150
        47919 => X"9E",  -- 158
        47920 => X"A3",  -- 163
        47921 => X"A9",  -- 169
        47922 => X"A0",  -- 160
        47923 => X"8D",  -- 141
        47924 => X"80",  -- 128
        47925 => X"7D",  -- 125
        47926 => X"8B",  -- 139
        47927 => X"A1",  -- 161
        47928 => X"AD",  -- 173
        47929 => X"A8",  -- 168
        47930 => X"AB",  -- 171
        47931 => X"B3",  -- 179
        47932 => X"A5",  -- 165
        47933 => X"A1",  -- 161
        47934 => X"B5",  -- 181
        47935 => X"B1",  -- 177
        47936 => X"B0",  -- 176
        47937 => X"B1",  -- 177
        47938 => X"A1",  -- 161
        47939 => X"A5",  -- 165
        47940 => X"A9",  -- 169
        47941 => X"A0",  -- 160
        47942 => X"A1",  -- 161
        47943 => X"A9",  -- 169
        47944 => X"9D",  -- 157
        47945 => X"AE",  -- 174
        47946 => X"A6",  -- 166
        47947 => X"AE",  -- 174
        47948 => X"B0",  -- 176
        47949 => X"B2",  -- 178
        47950 => X"C5",  -- 197
        47951 => X"BF",  -- 191
        47952 => X"B5",  -- 181
        47953 => X"B0",  -- 176
        47954 => X"AE",  -- 174
        47955 => X"B1",  -- 177
        47956 => X"B7",  -- 183
        47957 => X"BC",  -- 188
        47958 => X"C2",  -- 194
        47959 => X"C6",  -- 198
        47960 => X"BE",  -- 190
        47961 => X"BC",  -- 188
        47962 => X"BC",  -- 188
        47963 => X"BC",  -- 188
        47964 => X"C0",  -- 192
        47965 => X"C2",  -- 194
        47966 => X"C3",  -- 195
        47967 => X"C3",  -- 195
        47968 => X"C1",  -- 193
        47969 => X"C7",  -- 199
        47970 => X"CB",  -- 203
        47971 => X"CD",  -- 205
        47972 => X"CA",  -- 202
        47973 => X"C6",  -- 198
        47974 => X"C3",  -- 195
        47975 => X"C2",  -- 194
        47976 => X"B9",  -- 185
        47977 => X"B0",  -- 176
        47978 => X"A2",  -- 162
        47979 => X"9E",  -- 158
        47980 => X"AA",  -- 170
        47981 => X"B4",  -- 180
        47982 => X"A5",  -- 165
        47983 => X"8D",  -- 141
        47984 => X"86",  -- 134
        47985 => X"71",  -- 113
        47986 => X"51",  -- 81
        47987 => X"2C",  -- 44
        47988 => X"25",  -- 37
        47989 => X"35",  -- 53
        47990 => X"3C",  -- 60
        47991 => X"3C",  -- 60
        47992 => X"3A",  -- 58
        47993 => X"41",  -- 65
        47994 => X"48",  -- 72
        47995 => X"55",  -- 85
        47996 => X"65",  -- 101
        47997 => X"70",  -- 112
        47998 => X"7F",  -- 127
        47999 => X"95",  -- 149
        48000 => X"75",  -- 117
        48001 => X"71",  -- 113
        48002 => X"73",  -- 115
        48003 => X"7A",  -- 122
        48004 => X"7E",  -- 126
        48005 => X"7B",  -- 123
        48006 => X"78",  -- 120
        48007 => X"77",  -- 119
        48008 => X"76",  -- 118
        48009 => X"78",  -- 120
        48010 => X"75",  -- 117
        48011 => X"6E",  -- 110
        48012 => X"6B",  -- 107
        48013 => X"6E",  -- 110
        48014 => X"70",  -- 112
        48015 => X"70",  -- 112
        48016 => X"6F",  -- 111
        48017 => X"71",  -- 113
        48018 => X"72",  -- 114
        48019 => X"6F",  -- 111
        48020 => X"68",  -- 104
        48021 => X"5D",  -- 93
        48022 => X"55",  -- 85
        48023 => X"4F",  -- 79
        48024 => X"4D",  -- 77
        48025 => X"4B",  -- 75
        48026 => X"4A",  -- 74
        48027 => X"4B",  -- 75
        48028 => X"4A",  -- 74
        48029 => X"47",  -- 71
        48030 => X"46",  -- 70
        48031 => X"44",  -- 68
        48032 => X"4A",  -- 74
        48033 => X"4B",  -- 75
        48034 => X"66",  -- 102
        48035 => X"73",  -- 115
        48036 => X"5C",  -- 92
        48037 => X"55",  -- 85
        48038 => X"60",  -- 96
        48039 => X"60",  -- 96
        48040 => X"61",  -- 97
        48041 => X"6A",  -- 106
        48042 => X"65",  -- 101
        48043 => X"6E",  -- 110
        48044 => X"5C",  -- 92
        48045 => X"54",  -- 84
        48046 => X"60",  -- 96
        48047 => X"37",  -- 55
        48048 => X"11",  -- 17
        48049 => X"0A",  -- 10
        48050 => X"0B",  -- 11
        48051 => X"0F",  -- 15
        48052 => X"16",  -- 22
        48053 => X"28",  -- 40
        48054 => X"35",  -- 53
        48055 => X"32",  -- 50
        48056 => X"42",  -- 66
        48057 => X"59",  -- 89
        48058 => X"33",  -- 51
        48059 => X"35",  -- 53
        48060 => X"67",  -- 103
        48061 => X"32",  -- 50
        48062 => X"1D",  -- 29
        48063 => X"60",  -- 96
        48064 => X"59",  -- 89
        48065 => X"4C",  -- 76
        48066 => X"48",  -- 72
        48067 => X"4A",  -- 74
        48068 => X"47",  -- 71
        48069 => X"4C",  -- 76
        48070 => X"4B",  -- 75
        48071 => X"3E",  -- 62
        48072 => X"3D",  -- 61
        48073 => X"33",  -- 51
        48074 => X"2F",  -- 47
        48075 => X"33",  -- 51
        48076 => X"3D",  -- 61
        48077 => X"42",  -- 66
        48078 => X"43",  -- 67
        48079 => X"45",  -- 69
        48080 => X"56",  -- 86
        48081 => X"3D",  -- 61
        48082 => X"5B",  -- 91
        48083 => X"79",  -- 121
        48084 => X"65",  -- 101
        48085 => X"65",  -- 101
        48086 => X"79",  -- 121
        48087 => X"6C",  -- 108
        48088 => X"73",  -- 115
        48089 => X"7C",  -- 124
        48090 => X"82",  -- 130
        48091 => X"82",  -- 130
        48092 => X"85",  -- 133
        48093 => X"8A",  -- 138
        48094 => X"87",  -- 135
        48095 => X"80",  -- 128
        48096 => X"75",  -- 117
        48097 => X"7F",  -- 127
        48098 => X"81",  -- 129
        48099 => X"81",  -- 129
        48100 => X"85",  -- 133
        48101 => X"81",  -- 129
        48102 => X"78",  -- 120
        48103 => X"76",  -- 118
        48104 => X"71",  -- 113
        48105 => X"77",  -- 119
        48106 => X"85",  -- 133
        48107 => X"91",  -- 145
        48108 => X"8D",  -- 141
        48109 => X"79",  -- 121
        48110 => X"63",  -- 99
        48111 => X"56",  -- 86
        48112 => X"5F",  -- 95
        48113 => X"69",  -- 105
        48114 => X"64",  -- 100
        48115 => X"59",  -- 89
        48116 => X"5C",  -- 92
        48117 => X"63",  -- 99
        48118 => X"6C",  -- 108
        48119 => X"77",  -- 119
        48120 => X"69",  -- 105
        48121 => X"83",  -- 131
        48122 => X"76",  -- 118
        48123 => X"71",  -- 113
        48124 => X"85",  -- 133
        48125 => X"87",  -- 135
        48126 => X"95",  -- 149
        48127 => X"B2",  -- 178
        48128 => X"A1",  -- 161
        48129 => X"6F",  -- 111
        48130 => X"91",  -- 145
        48131 => X"D1",  -- 209
        48132 => X"E5",  -- 229
        48133 => X"DE",  -- 222
        48134 => X"C7",  -- 199
        48135 => X"BB",  -- 187
        48136 => X"90",  -- 144
        48137 => X"82",  -- 130
        48138 => X"7D",  -- 125
        48139 => X"6B",  -- 107
        48140 => X"3E",  -- 62
        48141 => X"0E",  -- 14
        48142 => X"01",  -- 1
        48143 => X"14",  -- 20
        48144 => X"0E",  -- 14
        48145 => X"0E",  -- 14
        48146 => X"07",  -- 7
        48147 => X"1F",  -- 31
        48148 => X"34",  -- 52
        48149 => X"35",  -- 53
        48150 => X"4D",  -- 77
        48151 => X"62",  -- 98
        48152 => X"74",  -- 116
        48153 => X"8B",  -- 139
        48154 => X"7D",  -- 125
        48155 => X"87",  -- 135
        48156 => X"8D",  -- 141
        48157 => X"79",  -- 121
        48158 => X"74",  -- 116
        48159 => X"90",  -- 144
        48160 => X"A2",  -- 162
        48161 => X"AC",  -- 172
        48162 => X"B2",  -- 178
        48163 => X"B9",  -- 185
        48164 => X"AA",  -- 170
        48165 => X"A2",  -- 162
        48166 => X"B8",  -- 184
        48167 => X"C0",  -- 192
        48168 => X"BD",  -- 189
        48169 => X"93",  -- 147
        48170 => X"93",  -- 147
        48171 => X"96",  -- 150
        48172 => X"69",  -- 105
        48173 => X"32",  -- 50
        48174 => X"32",  -- 50
        48175 => X"40",  -- 64
        48176 => X"3A",  -- 58
        48177 => X"3C",  -- 60
        48178 => X"3C",  -- 60
        48179 => X"3A",  -- 58
        48180 => X"36",  -- 54
        48181 => X"35",  -- 53
        48182 => X"38",  -- 56
        48183 => X"3C",  -- 60
        48184 => X"37",  -- 55
        48185 => X"37",  -- 55
        48186 => X"3C",  -- 60
        48187 => X"46",  -- 70
        48188 => X"4C",  -- 76
        48189 => X"48",  -- 72
        48190 => X"43",  -- 67
        48191 => X"3E",  -- 62
        48192 => X"3C",  -- 60
        48193 => X"38",  -- 56
        48194 => X"37",  -- 55
        48195 => X"38",  -- 56
        48196 => X"36",  -- 54
        48197 => X"33",  -- 51
        48198 => X"34",  -- 52
        48199 => X"38",  -- 56
        48200 => X"34",  -- 52
        48201 => X"35",  -- 53
        48202 => X"37",  -- 55
        48203 => X"37",  -- 55
        48204 => X"36",  -- 54
        48205 => X"36",  -- 54
        48206 => X"39",  -- 57
        48207 => X"3D",  -- 61
        48208 => X"3D",  -- 61
        48209 => X"3C",  -- 60
        48210 => X"39",  -- 57
        48211 => X"38",  -- 56
        48212 => X"3D",  -- 61
        48213 => X"44",  -- 68
        48214 => X"46",  -- 70
        48215 => X"42",  -- 66
        48216 => X"41",  -- 65
        48217 => X"44",  -- 68
        48218 => X"45",  -- 69
        48219 => X"43",  -- 67
        48220 => X"43",  -- 67
        48221 => X"45",  -- 69
        48222 => X"45",  -- 69
        48223 => X"43",  -- 67
        48224 => X"41",  -- 65
        48225 => X"46",  -- 70
        48226 => X"50",  -- 80
        48227 => X"6C",  -- 108
        48228 => X"87",  -- 135
        48229 => X"8C",  -- 140
        48230 => X"87",  -- 135
        48231 => X"8D",  -- 141
        48232 => X"90",  -- 144
        48233 => X"8C",  -- 140
        48234 => X"8D",  -- 141
        48235 => X"89",  -- 137
        48236 => X"94",  -- 148
        48237 => X"9D",  -- 157
        48238 => X"96",  -- 150
        48239 => X"9F",  -- 159
        48240 => X"A5",  -- 165
        48241 => X"AE",  -- 174
        48242 => X"AF",  -- 175
        48243 => X"A6",  -- 166
        48244 => X"8F",  -- 143
        48245 => X"77",  -- 119
        48246 => X"7D",  -- 125
        48247 => X"99",  -- 153
        48248 => X"AA",  -- 170
        48249 => X"9C",  -- 156
        48250 => X"B1",  -- 177
        48251 => X"B4",  -- 180
        48252 => X"A5",  -- 165
        48253 => X"AB",  -- 171
        48254 => X"AC",  -- 172
        48255 => X"A8",  -- 168
        48256 => X"AE",  -- 174
        48257 => X"AC",  -- 172
        48258 => X"A9",  -- 169
        48259 => X"A4",  -- 164
        48260 => X"A8",  -- 168
        48261 => X"A4",  -- 164
        48262 => X"9C",  -- 156
        48263 => X"AE",  -- 174
        48264 => X"A1",  -- 161
        48265 => X"AC",  -- 172
        48266 => X"AE",  -- 174
        48267 => X"AB",  -- 171
        48268 => X"AE",  -- 174
        48269 => X"B6",  -- 182
        48270 => X"C0",  -- 192
        48271 => X"C0",  -- 192
        48272 => X"B5",  -- 181
        48273 => X"B5",  -- 181
        48274 => X"B1",  -- 177
        48275 => X"AE",  -- 174
        48276 => X"B1",  -- 177
        48277 => X"BC",  -- 188
        48278 => X"C7",  -- 199
        48279 => X"CD",  -- 205
        48280 => X"BB",  -- 187
        48281 => X"BC",  -- 188
        48282 => X"BE",  -- 190
        48283 => X"BE",  -- 190
        48284 => X"C0",  -- 192
        48285 => X"C1",  -- 193
        48286 => X"C2",  -- 194
        48287 => X"C4",  -- 196
        48288 => X"C2",  -- 194
        48289 => X"C5",  -- 197
        48290 => X"C9",  -- 201
        48291 => X"CB",  -- 203
        48292 => X"CA",  -- 202
        48293 => X"C7",  -- 199
        48294 => X"C3",  -- 195
        48295 => X"C0",  -- 192
        48296 => X"B9",  -- 185
        48297 => X"B4",  -- 180
        48298 => X"A2",  -- 162
        48299 => X"91",  -- 145
        48300 => X"97",  -- 151
        48301 => X"A8",  -- 168
        48302 => X"A4",  -- 164
        48303 => X"8F",  -- 143
        48304 => X"70",  -- 112
        48305 => X"7B",  -- 123
        48306 => X"5A",  -- 90
        48307 => X"52",  -- 82
        48308 => X"3D",  -- 61
        48309 => X"22",  -- 34
        48310 => X"38",  -- 56
        48311 => X"2E",  -- 46
        48312 => X"34",  -- 52
        48313 => X"40",  -- 64
        48314 => X"4E",  -- 78
        48315 => X"5F",  -- 95
        48316 => X"6F",  -- 111
        48317 => X"73",  -- 115
        48318 => X"7C",  -- 124
        48319 => X"8F",  -- 143
        48320 => X"7E",  -- 126
        48321 => X"73",  -- 115
        48322 => X"6B",  -- 107
        48323 => X"6D",  -- 109
        48324 => X"70",  -- 112
        48325 => X"6F",  -- 111
        48326 => X"6D",  -- 109
        48327 => X"6E",  -- 110
        48328 => X"6B",  -- 107
        48329 => X"6D",  -- 109
        48330 => X"6B",  -- 107
        48331 => X"66",  -- 102
        48332 => X"66",  -- 102
        48333 => X"6B",  -- 107
        48334 => X"6C",  -- 108
        48335 => X"6A",  -- 106
        48336 => X"66",  -- 102
        48337 => X"6A",  -- 106
        48338 => X"6F",  -- 111
        48339 => X"70",  -- 112
        48340 => X"69",  -- 105
        48341 => X"60",  -- 96
        48342 => X"57",  -- 87
        48343 => X"50",  -- 80
        48344 => X"50",  -- 80
        48345 => X"51",  -- 81
        48346 => X"53",  -- 83
        48347 => X"54",  -- 84
        48348 => X"53",  -- 83
        48349 => X"4F",  -- 79
        48350 => X"4B",  -- 75
        48351 => X"46",  -- 70
        48352 => X"4D",  -- 77
        48353 => X"49",  -- 73
        48354 => X"5F",  -- 95
        48355 => X"6A",  -- 106
        48356 => X"56",  -- 86
        48357 => X"54",  -- 84
        48358 => X"63",  -- 99
        48359 => X"5C",  -- 92
        48360 => X"5D",  -- 93
        48361 => X"6C",  -- 108
        48362 => X"69",  -- 105
        48363 => X"6D",  -- 109
        48364 => X"55",  -- 85
        48365 => X"4D",  -- 77
        48366 => X"63",  -- 99
        48367 => X"40",  -- 64
        48368 => X"22",  -- 34
        48369 => X"15",  -- 21
        48370 => X"0D",  -- 13
        48371 => X"06",  -- 6
        48372 => X"05",  -- 5
        48373 => X"19",  -- 25
        48374 => X"30",  -- 48
        48375 => X"36",  -- 54
        48376 => X"3F",  -- 63
        48377 => X"57",  -- 87
        48378 => X"36",  -- 54
        48379 => X"22",  -- 34
        48380 => X"41",  -- 65
        48381 => X"1F",  -- 31
        48382 => X"4A",  -- 74
        48383 => X"5C",  -- 92
        48384 => X"57",  -- 87
        48385 => X"54",  -- 84
        48386 => X"4A",  -- 74
        48387 => X"48",  -- 72
        48388 => X"4E",  -- 78
        48389 => X"4B",  -- 75
        48390 => X"3C",  -- 60
        48391 => X"33",  -- 51
        48392 => X"3E",  -- 62
        48393 => X"34",  -- 52
        48394 => X"30",  -- 48
        48395 => X"35",  -- 53
        48396 => X"3E",  -- 62
        48397 => X"42",  -- 66
        48398 => X"43",  -- 67
        48399 => X"46",  -- 70
        48400 => X"56",  -- 86
        48401 => X"4C",  -- 76
        48402 => X"53",  -- 83
        48403 => X"6B",  -- 107
        48404 => X"73",  -- 115
        48405 => X"67",  -- 103
        48406 => X"66",  -- 102
        48407 => X"71",  -- 113
        48408 => X"62",  -- 98
        48409 => X"73",  -- 115
        48410 => X"84",  -- 132
        48411 => X"8B",  -- 139
        48412 => X"8E",  -- 142
        48413 => X"8E",  -- 142
        48414 => X"85",  -- 133
        48415 => X"7A",  -- 122
        48416 => X"7B",  -- 123
        48417 => X"7F",  -- 127
        48418 => X"78",  -- 120
        48419 => X"72",  -- 114
        48420 => X"76",  -- 118
        48421 => X"78",  -- 120
        48422 => X"78",  -- 120
        48423 => X"7C",  -- 124
        48424 => X"67",  -- 103
        48425 => X"6D",  -- 109
        48426 => X"78",  -- 120
        48427 => X"81",  -- 129
        48428 => X"7C",  -- 124
        48429 => X"6C",  -- 108
        48430 => X"60",  -- 96
        48431 => X"5B",  -- 91
        48432 => X"5F",  -- 95
        48433 => X"67",  -- 103
        48434 => X"60",  -- 96
        48435 => X"55",  -- 85
        48436 => X"5D",  -- 93
        48437 => X"69",  -- 105
        48438 => X"6C",  -- 108
        48439 => X"6E",  -- 110
        48440 => X"6F",  -- 111
        48441 => X"7F",  -- 127
        48442 => X"73",  -- 115
        48443 => X"87",  -- 135
        48444 => X"89",  -- 137
        48445 => X"58",  -- 88
        48446 => X"5B",  -- 91
        48447 => X"85",  -- 133
        48448 => X"B8",  -- 184
        48449 => X"7E",  -- 126
        48450 => X"59",  -- 89
        48451 => X"AB",  -- 171
        48452 => X"DF",  -- 223
        48453 => X"DB",  -- 219
        48454 => X"D1",  -- 209
        48455 => X"92",  -- 146
        48456 => X"89",  -- 137
        48457 => X"7F",  -- 127
        48458 => X"76",  -- 118
        48459 => X"57",  -- 87
        48460 => X"30",  -- 48
        48461 => X"12",  -- 18
        48462 => X"04",  -- 4
        48463 => X"0A",  -- 10
        48464 => X"07",  -- 7
        48465 => X"0A",  -- 10
        48466 => X"0D",  -- 13
        48467 => X"1B",  -- 27
        48468 => X"39",  -- 57
        48469 => X"4D",  -- 77
        48470 => X"55",  -- 85
        48471 => X"5C",  -- 92
        48472 => X"6B",  -- 107
        48473 => X"8B",  -- 139
        48474 => X"7A",  -- 122
        48475 => X"8C",  -- 140
        48476 => X"94",  -- 148
        48477 => X"7F",  -- 127
        48478 => X"6D",  -- 109
        48479 => X"8C",  -- 140
        48480 => X"A3",  -- 163
        48481 => X"AD",  -- 173
        48482 => X"B4",  -- 180
        48483 => X"B8",  -- 184
        48484 => X"A6",  -- 166
        48485 => X"9C",  -- 156
        48486 => X"B4",  -- 180
        48487 => X"BE",  -- 190
        48488 => X"C4",  -- 196
        48489 => X"92",  -- 146
        48490 => X"7D",  -- 125
        48491 => X"75",  -- 117
        48492 => X"6C",  -- 108
        48493 => X"32",  -- 50
        48494 => X"27",  -- 39
        48495 => X"39",  -- 57
        48496 => X"37",  -- 55
        48497 => X"3A",  -- 58
        48498 => X"3B",  -- 59
        48499 => X"39",  -- 57
        48500 => X"35",  -- 53
        48501 => X"33",  -- 51
        48502 => X"36",  -- 54
        48503 => X"39",  -- 57
        48504 => X"34",  -- 52
        48505 => X"34",  -- 52
        48506 => X"3A",  -- 58
        48507 => X"46",  -- 70
        48508 => X"4C",  -- 76
        48509 => X"4A",  -- 74
        48510 => X"44",  -- 68
        48511 => X"41",  -- 65
        48512 => X"3C",  -- 60
        48513 => X"37",  -- 55
        48514 => X"37",  -- 55
        48515 => X"39",  -- 57
        48516 => X"37",  -- 55
        48517 => X"32",  -- 50
        48518 => X"33",  -- 51
        48519 => X"37",  -- 55
        48520 => X"34",  -- 52
        48521 => X"34",  -- 52
        48522 => X"35",  -- 53
        48523 => X"35",  -- 53
        48524 => X"33",  -- 51
        48525 => X"34",  -- 52
        48526 => X"38",  -- 56
        48527 => X"3D",  -- 61
        48528 => X"3D",  -- 61
        48529 => X"3C",  -- 60
        48530 => X"39",  -- 57
        48531 => X"36",  -- 54
        48532 => X"3B",  -- 59
        48533 => X"44",  -- 68
        48534 => X"47",  -- 71
        48535 => X"43",  -- 67
        48536 => X"41",  -- 65
        48537 => X"47",  -- 71
        48538 => X"46",  -- 70
        48539 => X"41",  -- 65
        48540 => X"41",  -- 65
        48541 => X"46",  -- 70
        48542 => X"48",  -- 72
        48543 => X"42",  -- 66
        48544 => X"46",  -- 70
        48545 => X"4C",  -- 76
        48546 => X"58",  -- 88
        48547 => X"74",  -- 116
        48548 => X"8D",  -- 141
        48549 => X"8F",  -- 143
        48550 => X"88",  -- 136
        48551 => X"8F",  -- 143
        48552 => X"8C",  -- 140
        48553 => X"87",  -- 135
        48554 => X"8A",  -- 138
        48555 => X"88",  -- 136
        48556 => X"97",  -- 151
        48557 => X"A3",  -- 163
        48558 => X"A1",  -- 161
        48559 => X"AB",  -- 171
        48560 => X"AD",  -- 173
        48561 => X"B2",  -- 178
        48562 => X"B3",  -- 179
        48563 => X"B0",  -- 176
        48564 => X"9E",  -- 158
        48565 => X"82",  -- 130
        48566 => X"79",  -- 121
        48567 => X"89",  -- 137
        48568 => X"9F",  -- 159
        48569 => X"8B",  -- 139
        48570 => X"B1",  -- 177
        48571 => X"B4",  -- 180
        48572 => X"A7",  -- 167
        48573 => X"B1",  -- 177
        48574 => X"A6",  -- 166
        48575 => X"A1",  -- 161
        48576 => X"AB",  -- 171
        48577 => X"A9",  -- 169
        48578 => X"AF",  -- 175
        48579 => X"A5",  -- 165
        48580 => X"A8",  -- 168
        48581 => X"A6",  -- 166
        48582 => X"96",  -- 150
        48583 => X"B1",  -- 177
        48584 => X"A5",  -- 165
        48585 => X"AA",  -- 170
        48586 => X"B5",  -- 181
        48587 => X"AB",  -- 171
        48588 => X"AB",  -- 171
        48589 => X"B9",  -- 185
        48590 => X"BB",  -- 187
        48591 => X"C2",  -- 194
        48592 => X"B9",  -- 185
        48593 => X"BD",  -- 189
        48594 => X"B8",  -- 184
        48595 => X"AF",  -- 175
        48596 => X"AD",  -- 173
        48597 => X"B9",  -- 185
        48598 => X"C9",  -- 201
        48599 => X"D0",  -- 208
        48600 => X"BA",  -- 186
        48601 => X"BC",  -- 188
        48602 => X"C0",  -- 192
        48603 => X"C0",  -- 192
        48604 => X"BF",  -- 191
        48605 => X"C0",  -- 192
        48606 => X"C3",  -- 195
        48607 => X"C6",  -- 198
        48608 => X"C3",  -- 195
        48609 => X"C4",  -- 196
        48610 => X"C7",  -- 199
        48611 => X"CA",  -- 202
        48612 => X"CB",  -- 203
        48613 => X"C8",  -- 200
        48614 => X"C3",  -- 195
        48615 => X"BF",  -- 191
        48616 => X"B7",  -- 183
        48617 => X"B8",  -- 184
        48618 => X"A3",  -- 163
        48619 => X"86",  -- 134
        48620 => X"84",  -- 132
        48621 => X"98",  -- 152
        48622 => X"9C",  -- 156
        48623 => X"8D",  -- 141
        48624 => X"67",  -- 103
        48625 => X"75",  -- 117
        48626 => X"77",  -- 119
        48627 => X"43",  -- 67
        48628 => X"25",  -- 37
        48629 => X"31",  -- 49
        48630 => X"30",  -- 48
        48631 => X"35",  -- 53
        48632 => X"2A",  -- 42
        48633 => X"3A",  -- 58
        48634 => X"4F",  -- 79
        48635 => X"67",  -- 103
        48636 => X"78",  -- 120
        48637 => X"79",  -- 121
        48638 => X"7D",  -- 125
        48639 => X"8C",  -- 140
        48640 => X"6E",  -- 110
        48641 => X"6B",  -- 107
        48642 => X"69",  -- 105
        48643 => X"69",  -- 105
        48644 => X"6B",  -- 107
        48645 => X"6B",  -- 107
        48646 => X"69",  -- 105
        48647 => X"67",  -- 103
        48648 => X"61",  -- 97
        48649 => X"5E",  -- 94
        48650 => X"5C",  -- 92
        48651 => X"5B",  -- 91
        48652 => X"5D",  -- 93
        48653 => X"5F",  -- 95
        48654 => X"5F",  -- 95
        48655 => X"5E",  -- 94
        48656 => X"5F",  -- 95
        48657 => X"60",  -- 96
        48658 => X"61",  -- 97
        48659 => X"62",  -- 98
        48660 => X"62",  -- 98
        48661 => X"5B",  -- 91
        48662 => X"52",  -- 82
        48663 => X"4B",  -- 75
        48664 => X"4A",  -- 74
        48665 => X"4C",  -- 76
        48666 => X"4E",  -- 78
        48667 => X"53",  -- 83
        48668 => X"56",  -- 86
        48669 => X"54",  -- 84
        48670 => X"51",  -- 81
        48671 => X"4C",  -- 76
        48672 => X"4C",  -- 76
        48673 => X"4B",  -- 75
        48674 => X"58",  -- 88
        48675 => X"5D",  -- 93
        48676 => X"55",  -- 85
        48677 => X"5B",  -- 91
        48678 => X"60",  -- 96
        48679 => X"55",  -- 85
        48680 => X"58",  -- 88
        48681 => X"6E",  -- 110
        48682 => X"6E",  -- 110
        48683 => X"66",  -- 102
        48684 => X"54",  -- 84
        48685 => X"58",  -- 88
        48686 => X"65",  -- 101
        48687 => X"43",  -- 67
        48688 => X"2F",  -- 47
        48689 => X"1F",  -- 31
        48690 => X"1D",  -- 29
        48691 => X"0C",  -- 12
        48692 => X"17",  -- 23
        48693 => X"17",  -- 23
        48694 => X"24",  -- 36
        48695 => X"3C",  -- 60
        48696 => X"4C",  -- 76
        48697 => X"4E",  -- 78
        48698 => X"23",  -- 35
        48699 => X"3A",  -- 58
        48700 => X"2B",  -- 43
        48701 => X"2E",  -- 46
        48702 => X"5C",  -- 92
        48703 => X"63",  -- 99
        48704 => X"55",  -- 85
        48705 => X"54",  -- 84
        48706 => X"4A",  -- 74
        48707 => X"3D",  -- 61
        48708 => X"48",  -- 72
        48709 => X"3F",  -- 63
        48710 => X"31",  -- 49
        48711 => X"4A",  -- 74
        48712 => X"39",  -- 57
        48713 => X"2C",  -- 44
        48714 => X"2C",  -- 44
        48715 => X"33",  -- 51
        48716 => X"35",  -- 53
        48717 => X"39",  -- 57
        48718 => X"42",  -- 66
        48719 => X"45",  -- 69
        48720 => X"48",  -- 72
        48721 => X"53",  -- 83
        48722 => X"60",  -- 96
        48723 => X"68",  -- 104
        48724 => X"65",  -- 101
        48725 => X"78",  -- 120
        48726 => X"6E",  -- 110
        48727 => X"76",  -- 118
        48728 => X"71",  -- 113
        48729 => X"72",  -- 114
        48730 => X"76",  -- 118
        48731 => X"86",  -- 134
        48732 => X"8F",  -- 143
        48733 => X"84",  -- 132
        48734 => X"7E",  -- 126
        48735 => X"89",  -- 137
        48736 => X"83",  -- 131
        48737 => X"7E",  -- 126
        48738 => X"87",  -- 135
        48739 => X"70",  -- 112
        48740 => X"82",  -- 130
        48741 => X"77",  -- 119
        48742 => X"84",  -- 132
        48743 => X"7A",  -- 122
        48744 => X"75",  -- 117
        48745 => X"79",  -- 121
        48746 => X"67",  -- 103
        48747 => X"74",  -- 116
        48748 => X"7D",  -- 125
        48749 => X"6E",  -- 110
        48750 => X"69",  -- 105
        48751 => X"5A",  -- 90
        48752 => X"5B",  -- 91
        48753 => X"6B",  -- 107
        48754 => X"73",  -- 115
        48755 => X"69",  -- 105
        48756 => X"61",  -- 97
        48757 => X"65",  -- 101
        48758 => X"6C",  -- 108
        48759 => X"6E",  -- 110
        48760 => X"65",  -- 101
        48761 => X"7D",  -- 125
        48762 => X"7A",  -- 122
        48763 => X"81",  -- 129
        48764 => X"85",  -- 133
        48765 => X"40",  -- 64
        48766 => X"12",  -- 18
        48767 => X"36",  -- 54
        48768 => X"7B",  -- 123
        48769 => X"A8",  -- 168
        48770 => X"58",  -- 88
        48771 => X"64",  -- 100
        48772 => X"D8",  -- 216
        48773 => X"DC",  -- 220
        48774 => X"CD",  -- 205
        48775 => X"9E",  -- 158
        48776 => X"93",  -- 147
        48777 => X"91",  -- 145
        48778 => X"6C",  -- 108
        48779 => X"4C",  -- 76
        48780 => X"25",  -- 37
        48781 => X"06",  -- 6
        48782 => X"0C",  -- 12
        48783 => X"01",  -- 1
        48784 => X"09",  -- 9
        48785 => X"07",  -- 7
        48786 => X"1C",  -- 28
        48787 => X"22",  -- 34
        48788 => X"43",  -- 67
        48789 => X"67",  -- 103
        48790 => X"62",  -- 98
        48791 => X"5D",  -- 93
        48792 => X"67",  -- 103
        48793 => X"85",  -- 133
        48794 => X"8C",  -- 140
        48795 => X"84",  -- 132
        48796 => X"97",  -- 151
        48797 => X"9C",  -- 156
        48798 => X"67",  -- 103
        48799 => X"88",  -- 136
        48800 => X"8F",  -- 143
        48801 => X"BA",  -- 186
        48802 => X"B2",  -- 178
        48803 => X"B4",  -- 180
        48804 => X"B2",  -- 178
        48805 => X"93",  -- 147
        48806 => X"A7",  -- 167
        48807 => X"B8",  -- 184
        48808 => X"C4",  -- 196
        48809 => X"9D",  -- 157
        48810 => X"6B",  -- 107
        48811 => X"5D",  -- 93
        48812 => X"54",  -- 84
        48813 => X"33",  -- 51
        48814 => X"29",  -- 41
        48815 => X"2B",  -- 43
        48816 => X"31",  -- 49
        48817 => X"36",  -- 54
        48818 => X"38",  -- 56
        48819 => X"34",  -- 52
        48820 => X"30",  -- 48
        48821 => X"31",  -- 49
        48822 => X"34",  -- 52
        48823 => X"35",  -- 53
        48824 => X"39",  -- 57
        48825 => X"2E",  -- 46
        48826 => X"2D",  -- 45
        48827 => X"3E",  -- 62
        48828 => X"4C",  -- 76
        48829 => X"4C",  -- 76
        48830 => X"43",  -- 67
        48831 => X"3E",  -- 62
        48832 => X"3F",  -- 63
        48833 => X"3A",  -- 58
        48834 => X"39",  -- 57
        48835 => X"3A",  -- 58
        48836 => X"38",  -- 56
        48837 => X"34",  -- 52
        48838 => X"35",  -- 53
        48839 => X"3A",  -- 58
        48840 => X"35",  -- 53
        48841 => X"31",  -- 49
        48842 => X"30",  -- 48
        48843 => X"33",  -- 51
        48844 => X"35",  -- 53
        48845 => X"36",  -- 54
        48846 => X"38",  -- 56
        48847 => X"3C",  -- 60
        48848 => X"3B",  -- 59
        48849 => X"3D",  -- 61
        48850 => X"3C",  -- 60
        48851 => X"39",  -- 57
        48852 => X"39",  -- 57
        48853 => X"3D",  -- 61
        48854 => X"43",  -- 67
        48855 => X"42",  -- 66
        48856 => X"43",  -- 67
        48857 => X"45",  -- 69
        48858 => X"46",  -- 70
        48859 => X"41",  -- 65
        48860 => X"3C",  -- 60
        48861 => X"44",  -- 68
        48862 => X"49",  -- 73
        48863 => X"40",  -- 64
        48864 => X"4C",  -- 76
        48865 => X"43",  -- 67
        48866 => X"5D",  -- 93
        48867 => X"81",  -- 129
        48868 => X"8A",  -- 138
        48869 => X"8A",  -- 138
        48870 => X"8D",  -- 141
        48871 => X"89",  -- 137
        48872 => X"85",  -- 133
        48873 => X"80",  -- 128
        48874 => X"82",  -- 130
        48875 => X"8F",  -- 143
        48876 => X"99",  -- 153
        48877 => X"9E",  -- 158
        48878 => X"A4",  -- 164
        48879 => X"AA",  -- 170
        48880 => X"AE",  -- 174
        48881 => X"AE",  -- 174
        48882 => X"B3",  -- 179
        48883 => X"AD",  -- 173
        48884 => X"B3",  -- 179
        48885 => X"96",  -- 150
        48886 => X"87",  -- 135
        48887 => X"84",  -- 132
        48888 => X"87",  -- 135
        48889 => X"97",  -- 151
        48890 => X"93",  -- 147
        48891 => X"9B",  -- 155
        48892 => X"A5",  -- 165
        48893 => X"A2",  -- 162
        48894 => X"A6",  -- 166
        48895 => X"A3",  -- 163
        48896 => X"A2",  -- 162
        48897 => X"A5",  -- 165
        48898 => X"A8",  -- 168
        48899 => X"A9",  -- 169
        48900 => X"AB",  -- 171
        48901 => X"AC",  -- 172
        48902 => X"A9",  -- 169
        48903 => X"A5",  -- 165
        48904 => X"AD",  -- 173
        48905 => X"AC",  -- 172
        48906 => X"AB",  -- 171
        48907 => X"AB",  -- 171
        48908 => X"B3",  -- 179
        48909 => X"C0",  -- 192
        48910 => X"C2",  -- 194
        48911 => X"BF",  -- 191
        48912 => X"BB",  -- 187
        48913 => X"BC",  -- 188
        48914 => X"B9",  -- 185
        48915 => X"B1",  -- 177
        48916 => X"B5",  -- 181
        48917 => X"C1",  -- 193
        48918 => X"C8",  -- 200
        48919 => X"C6",  -- 198
        48920 => X"BA",  -- 186
        48921 => X"B9",  -- 185
        48922 => X"BE",  -- 190
        48923 => X"C3",  -- 195
        48924 => X"C3",  -- 195
        48925 => X"BF",  -- 191
        48926 => X"C2",  -- 194
        48927 => X"C7",  -- 199
        48928 => X"C7",  -- 199
        48929 => X"C4",  -- 196
        48930 => X"C5",  -- 197
        48931 => X"CB",  -- 203
        48932 => X"CD",  -- 205
        48933 => X"C8",  -- 200
        48934 => X"C3",  -- 195
        48935 => X"C1",  -- 193
        48936 => X"AB",  -- 171
        48937 => X"AF",  -- 175
        48938 => X"B1",  -- 177
        48939 => X"9F",  -- 159
        48940 => X"80",  -- 128
        48941 => X"78",  -- 120
        48942 => X"87",  -- 135
        48943 => X"92",  -- 146
        48944 => X"7A",  -- 122
        48945 => X"62",  -- 98
        48946 => X"5E",  -- 94
        48947 => X"5D",  -- 93
        48948 => X"42",  -- 66
        48949 => X"2B",  -- 43
        48950 => X"2B",  -- 43
        48951 => X"2A",  -- 42
        48952 => X"3D",  -- 61
        48953 => X"3A",  -- 58
        48954 => X"4A",  -- 74
        48955 => X"67",  -- 103
        48956 => X"7C",  -- 124
        48957 => X"82",  -- 130
        48958 => X"87",  -- 135
        48959 => X"8E",  -- 142
        48960 => X"5D",  -- 93
        48961 => X"5D",  -- 93
        48962 => X"5D",  -- 93
        48963 => X"5D",  -- 93
        48964 => X"5E",  -- 94
        48965 => X"5C",  -- 92
        48966 => X"5A",  -- 90
        48967 => X"58",  -- 88
        48968 => X"56",  -- 86
        48969 => X"55",  -- 85
        48970 => X"53",  -- 83
        48971 => X"53",  -- 83
        48972 => X"54",  -- 84
        48973 => X"55",  -- 85
        48974 => X"56",  -- 86
        48975 => X"56",  -- 86
        48976 => X"57",  -- 87
        48977 => X"5A",  -- 90
        48978 => X"5C",  -- 92
        48979 => X"5A",  -- 90
        48980 => X"55",  -- 85
        48981 => X"50",  -- 80
        48982 => X"4F",  -- 79
        48983 => X"4F",  -- 79
        48984 => X"4F",  -- 79
        48985 => X"4D",  -- 77
        48986 => X"4C",  -- 76
        48987 => X"4D",  -- 77
        48988 => X"4E",  -- 78
        48989 => X"4F",  -- 79
        48990 => X"4B",  -- 75
        48991 => X"48",  -- 72
        48992 => X"48",  -- 72
        48993 => X"47",  -- 71
        48994 => X"51",  -- 81
        48995 => X"56",  -- 86
        48996 => X"53",  -- 83
        48997 => X"5C",  -- 92
        48998 => X"62",  -- 98
        48999 => X"57",  -- 87
        49000 => X"59",  -- 89
        49001 => X"6F",  -- 111
        49002 => X"6F",  -- 111
        49003 => X"61",  -- 97
        49004 => X"4F",  -- 79
        49005 => X"56",  -- 86
        49006 => X"64",  -- 100
        49007 => X"46",  -- 70
        49008 => X"3F",  -- 63
        49009 => X"30",  -- 48
        49010 => X"28",  -- 40
        49011 => X"0F",  -- 15
        49012 => X"13",  -- 19
        49013 => X"0F",  -- 15
        49014 => X"13",  -- 19
        49015 => X"23",  -- 35
        49016 => X"39",  -- 57
        49017 => X"41",  -- 65
        49018 => X"3C",  -- 60
        49019 => X"32",  -- 50
        49020 => X"2E",  -- 46
        49021 => X"4F",  -- 79
        49022 => X"67",  -- 103
        49023 => X"67",  -- 103
        49024 => X"51",  -- 81
        49025 => X"4E",  -- 78
        49026 => X"44",  -- 68
        49027 => X"3C",  -- 60
        49028 => X"4B",  -- 75
        49029 => X"46",  -- 70
        49030 => X"37",  -- 55
        49031 => X"4C",  -- 76
        49032 => X"4B",  -- 75
        49033 => X"32",  -- 50
        49034 => X"25",  -- 37
        49035 => X"2A",  -- 42
        49036 => X"36",  -- 54
        49037 => X"3F",  -- 63
        49038 => X"43",  -- 67
        49039 => X"40",  -- 64
        49040 => X"4A",  -- 74
        49041 => X"57",  -- 87
        49042 => X"67",  -- 103
        49043 => X"70",  -- 112
        49044 => X"6A",  -- 106
        49045 => X"78",  -- 120
        49046 => X"6B",  -- 107
        49047 => X"71",  -- 113
        49048 => X"6B",  -- 107
        49049 => X"73",  -- 115
        49050 => X"7C",  -- 124
        49051 => X"86",  -- 134
        49052 => X"87",  -- 135
        49053 => X"77",  -- 119
        49054 => X"74",  -- 116
        49055 => X"83",  -- 131
        49056 => X"7F",  -- 127
        49057 => X"80",  -- 128
        49058 => X"81",  -- 129
        49059 => X"7D",  -- 125
        49060 => X"8A",  -- 138
        49061 => X"85",  -- 133
        49062 => X"85",  -- 133
        49063 => X"86",  -- 134
        49064 => X"7B",  -- 123
        49065 => X"7E",  -- 126
        49066 => X"65",  -- 101
        49067 => X"67",  -- 103
        49068 => X"75",  -- 117
        49069 => X"75",  -- 117
        49070 => X"68",  -- 104
        49071 => X"46",  -- 70
        49072 => X"60",  -- 96
        49073 => X"67",  -- 103
        49074 => X"6E",  -- 110
        49075 => X"70",  -- 112
        49076 => X"6F",  -- 111
        49077 => X"70",  -- 112
        49078 => X"71",  -- 113
        49079 => X"74",  -- 116
        49080 => X"7E",  -- 126
        49081 => X"7B",  -- 123
        49082 => X"71",  -- 113
        49083 => X"78",  -- 120
        49084 => X"8D",  -- 141
        49085 => X"77",  -- 119
        49086 => X"3A",  -- 58
        49087 => X"0E",  -- 14
        49088 => X"2E",  -- 46
        49089 => X"99",  -- 153
        49090 => X"8F",  -- 143
        49091 => X"65",  -- 101
        49092 => X"C0",  -- 192
        49093 => X"DC",  -- 220
        49094 => X"C1",  -- 193
        49095 => X"90",  -- 144
        49096 => X"96",  -- 150
        49097 => X"94",  -- 148
        49098 => X"78",  -- 120
        49099 => X"48",  -- 72
        49100 => X"16",  -- 22
        49101 => X"05",  -- 5
        49102 => X"0D",  -- 13
        49103 => X"03",  -- 3
        49104 => X"0F",  -- 15
        49105 => X"10",  -- 16
        49106 => X"23",  -- 35
        49107 => X"2B",  -- 43
        49108 => X"4A",  -- 74
        49109 => X"6E",  -- 110
        49110 => X"6B",  -- 107
        49111 => X"67",  -- 103
        49112 => X"61",  -- 97
        49113 => X"7F",  -- 127
        49114 => X"8B",  -- 139
        49115 => X"8C",  -- 140
        49116 => X"92",  -- 146
        49117 => X"9D",  -- 157
        49118 => X"6C",  -- 108
        49119 => X"83",  -- 131
        49120 => X"8C",  -- 140
        49121 => X"B5",  -- 181
        49122 => X"AD",  -- 173
        49123 => X"B1",  -- 177
        49124 => X"AD",  -- 173
        49125 => X"93",  -- 147
        49126 => X"A3",  -- 163
        49127 => X"B2",  -- 178
        49128 => X"BE",  -- 190
        49129 => X"91",  -- 145
        49130 => X"5E",  -- 94
        49131 => X"4F",  -- 79
        49132 => X"4C",  -- 76
        49133 => X"25",  -- 37
        49134 => X"26",  -- 38
        49135 => X"34",  -- 52
        49136 => X"31",  -- 49
        49137 => X"36",  -- 54
        49138 => X"37",  -- 55
        49139 => X"32",  -- 50
        49140 => X"2F",  -- 47
        49141 => X"30",  -- 48
        49142 => X"33",  -- 51
        49143 => X"34",  -- 52
        49144 => X"36",  -- 54
        49145 => X"2C",  -- 44
        49146 => X"2D",  -- 45
        49147 => X"3D",  -- 61
        49148 => X"4C",  -- 76
        49149 => X"4C",  -- 76
        49150 => X"45",  -- 69
        49151 => X"40",  -- 64
        49152 => X"3F",  -- 63
        49153 => X"3B",  -- 59
        49154 => X"3A",  -- 58
        49155 => X"3B",  -- 59
        49156 => X"39",  -- 57
        49157 => X"35",  -- 53
        49158 => X"36",  -- 54
        49159 => X"39",  -- 57
        49160 => X"35",  -- 53
        49161 => X"30",  -- 48
        49162 => X"2E",  -- 46
        49163 => X"31",  -- 49
        49164 => X"35",  -- 53
        49165 => X"36",  -- 54
        49166 => X"38",  -- 56
        49167 => X"3B",  -- 59
        49168 => X"39",  -- 57
        49169 => X"39",  -- 57
        49170 => X"39",  -- 57
        49171 => X"37",  -- 55
        49172 => X"3B",  -- 59
        49173 => X"43",  -- 67
        49174 => X"47",  -- 71
        49175 => X"48",  -- 72
        49176 => X"47",  -- 71
        49177 => X"46",  -- 70
        49178 => X"49",  -- 73
        49179 => X"47",  -- 71
        49180 => X"42",  -- 66
        49181 => X"45",  -- 69
        49182 => X"49",  -- 73
        49183 => X"45",  -- 69
        49184 => X"47",  -- 71
        49185 => X"59",  -- 89
        49186 => X"77",  -- 119
        49187 => X"8F",  -- 143
        49188 => X"95",  -- 149
        49189 => X"93",  -- 147
        49190 => X"91",  -- 145
        49191 => X"8B",  -- 139
        49192 => X"88",  -- 136
        49193 => X"85",  -- 133
        49194 => X"87",  -- 135
        49195 => X"8D",  -- 141
        49196 => X"93",  -- 147
        49197 => X"99",  -- 153
        49198 => X"9E",  -- 158
        49199 => X"A3",  -- 163
        49200 => X"A3",  -- 163
        49201 => X"9E",  -- 158
        49202 => X"A8",  -- 168
        49203 => X"B0",  -- 176
        49204 => X"BA",  -- 186
        49205 => X"9F",  -- 159
        49206 => X"92",  -- 146
        49207 => X"8D",  -- 141
        49208 => X"8B",  -- 139
        49209 => X"94",  -- 148
        49210 => X"93",  -- 147
        49211 => X"9B",  -- 155
        49212 => X"9D",  -- 157
        49213 => X"A0",  -- 160
        49214 => X"A8",  -- 168
        49215 => X"A0",  -- 160
        49216 => X"A0",  -- 160
        49217 => X"A0",  -- 160
        49218 => X"A4",  -- 164
        49219 => X"A7",  -- 167
        49220 => X"AA",  -- 170
        49221 => X"A8",  -- 168
        49222 => X"A6",  -- 166
        49223 => X"A4",  -- 164
        49224 => X"B0",  -- 176
        49225 => X"AF",  -- 175
        49226 => X"AF",  -- 175
        49227 => X"B2",  -- 178
        49228 => X"B6",  -- 182
        49229 => X"BA",  -- 186
        49230 => X"BD",  -- 189
        49231 => X"BF",  -- 191
        49232 => X"BA",  -- 186
        49233 => X"BC",  -- 188
        49234 => X"B8",  -- 184
        49235 => X"B1",  -- 177
        49236 => X"B3",  -- 179
        49237 => X"BF",  -- 191
        49238 => X"C4",  -- 196
        49239 => X"C3",  -- 195
        49240 => X"B7",  -- 183
        49241 => X"B7",  -- 183
        49242 => X"BA",  -- 186
        49243 => X"C0",  -- 192
        49244 => X"C2",  -- 194
        49245 => X"C0",  -- 192
        49246 => X"C2",  -- 194
        49247 => X"C7",  -- 199
        49248 => X"C6",  -- 198
        49249 => X"C3",  -- 195
        49250 => X"C3",  -- 195
        49251 => X"C8",  -- 200
        49252 => X"CA",  -- 202
        49253 => X"C6",  -- 198
        49254 => X"C2",  -- 194
        49255 => X"C0",  -- 192
        49256 => X"C2",  -- 194
        49257 => X"A2",  -- 162
        49258 => X"9E",  -- 158
        49259 => X"AC",  -- 172
        49260 => X"96",  -- 150
        49261 => X"70",  -- 112
        49262 => X"6C",  -- 108
        49263 => X"80",  -- 128
        49264 => X"7F",  -- 127
        49265 => X"64",  -- 100
        49266 => X"51",  -- 81
        49267 => X"4E",  -- 78
        49268 => X"46",  -- 70
        49269 => X"3C",  -- 60
        49270 => X"34",  -- 52
        49271 => X"2F",  -- 47
        49272 => X"44",  -- 68
        49273 => X"48",  -- 72
        49274 => X"54",  -- 84
        49275 => X"65",  -- 101
        49276 => X"75",  -- 117
        49277 => X"85",  -- 133
        49278 => X"93",  -- 147
        49279 => X"9C",  -- 156
        49280 => X"47",  -- 71
        49281 => X"49",  -- 73
        49282 => X"4C",  -- 76
        49283 => X"4C",  -- 76
        49284 => X"4A",  -- 74
        49285 => X"48",  -- 72
        49286 => X"46",  -- 70
        49287 => X"45",  -- 69
        49288 => X"4A",  -- 74
        49289 => X"4B",  -- 75
        49290 => X"4C",  -- 76
        49291 => X"4C",  -- 76
        49292 => X"4B",  -- 75
        49293 => X"4C",  -- 76
        49294 => X"4D",  -- 77
        49295 => X"50",  -- 80
        49296 => X"4F",  -- 79
        49297 => X"53",  -- 83
        49298 => X"56",  -- 86
        49299 => X"50",  -- 80
        49300 => X"49",  -- 73
        49301 => X"46",  -- 70
        49302 => X"4A",  -- 74
        49303 => X"51",  -- 81
        49304 => X"4F",  -- 79
        49305 => X"4C",  -- 76
        49306 => X"47",  -- 71
        49307 => X"46",  -- 70
        49308 => X"46",  -- 70
        49309 => X"46",  -- 70
        49310 => X"44",  -- 68
        49311 => X"41",  -- 65
        49312 => X"3F",  -- 63
        49313 => X"3E",  -- 62
        49314 => X"44",  -- 68
        49315 => X"49",  -- 73
        49316 => X"4C",  -- 76
        49317 => X"53",  -- 83
        49318 => X"58",  -- 88
        49319 => X"50",  -- 80
        49320 => X"56",  -- 86
        49321 => X"6D",  -- 109
        49322 => X"6B",  -- 107
        49323 => X"57",  -- 87
        49324 => X"4A",  -- 74
        49325 => X"57",  -- 87
        49326 => X"63",  -- 99
        49327 => X"48",  -- 72
        49328 => X"48",  -- 72
        49329 => X"3D",  -- 61
        49330 => X"35",  -- 53
        49331 => X"15",  -- 21
        49332 => X"18",  -- 24
        49333 => X"13",  -- 19
        49334 => X"10",  -- 16
        49335 => X"15",  -- 21
        49336 => X"23",  -- 35
        49337 => X"33",  -- 51
        49338 => X"54",  -- 84
        49339 => X"30",  -- 48
        49340 => X"38",  -- 56
        49341 => X"6C",  -- 108
        49342 => X"6D",  -- 109
        49343 => X"62",  -- 98
        49344 => X"53",  -- 83
        49345 => X"4D",  -- 77
        49346 => X"44",  -- 68
        49347 => X"3D",  -- 61
        49348 => X"49",  -- 73
        49349 => X"45",  -- 69
        49350 => X"34",  -- 52
        49351 => X"3F",  -- 63
        49352 => X"4F",  -- 79
        49353 => X"35",  -- 53
        49354 => X"22",  -- 34
        49355 => X"27",  -- 39
        49356 => X"37",  -- 55
        49357 => X"40",  -- 64
        49358 => X"3F",  -- 63
        49359 => X"3C",  -- 60
        49360 => X"4C",  -- 76
        49361 => X"59",  -- 89
        49362 => X"69",  -- 105
        49363 => X"72",  -- 114
        49364 => X"6A",  -- 106
        49365 => X"76",  -- 118
        49366 => X"6A",  -- 106
        49367 => X"73",  -- 115
        49368 => X"77",  -- 119
        49369 => X"7E",  -- 126
        49370 => X"83",  -- 131
        49371 => X"8C",  -- 140
        49372 => X"8D",  -- 141
        49373 => X"7F",  -- 127
        49374 => X"7A",  -- 122
        49375 => X"84",  -- 132
        49376 => X"7A",  -- 122
        49377 => X"82",  -- 130
        49378 => X"7B",  -- 123
        49379 => X"81",  -- 129
        49380 => X"87",  -- 135
        49381 => X"85",  -- 133
        49382 => X"7A",  -- 122
        49383 => X"87",  -- 135
        49384 => X"88",  -- 136
        49385 => X"83",  -- 131
        49386 => X"6F",  -- 111
        49387 => X"6F",  -- 111
        49388 => X"78",  -- 120
        49389 => X"75",  -- 117
        49390 => X"67",  -- 103
        49391 => X"4B",  -- 75
        49392 => X"58",  -- 88
        49393 => X"57",  -- 87
        49394 => X"5E",  -- 94
        49395 => X"6D",  -- 109
        49396 => X"75",  -- 117
        49397 => X"77",  -- 119
        49398 => X"76",  -- 118
        49399 => X"77",  -- 119
        49400 => X"7D",  -- 125
        49401 => X"74",  -- 116
        49402 => X"79",  -- 121
        49403 => X"82",  -- 130
        49404 => X"89",  -- 137
        49405 => X"93",  -- 147
        49406 => X"73",  -- 115
        49407 => X"31",  -- 49
        49408 => X"2C",  -- 44
        49409 => X"97",  -- 151
        49410 => X"C6",  -- 198
        49411 => X"69",  -- 105
        49412 => X"A0",  -- 160
        49413 => X"D2",  -- 210
        49414 => X"AF",  -- 175
        49415 => X"8D",  -- 141
        49416 => X"88",  -- 136
        49417 => X"82",  -- 130
        49418 => X"7C",  -- 124
        49419 => X"45",  -- 69
        49420 => X"08",  -- 8
        49421 => X"04",  -- 4
        49422 => X"0B",  -- 11
        49423 => X"03",  -- 3
        49424 => X"12",  -- 18
        49425 => X"1A",  -- 26
        49426 => X"2C",  -- 44
        49427 => X"3C",  -- 60
        49428 => X"53",  -- 83
        49429 => X"71",  -- 113
        49430 => X"6C",  -- 108
        49431 => X"67",  -- 103
        49432 => X"60",  -- 96
        49433 => X"7C",  -- 124
        49434 => X"8E",  -- 142
        49435 => X"9B",  -- 155
        49436 => X"8E",  -- 142
        49437 => X"A0",  -- 160
        49438 => X"77",  -- 119
        49439 => X"81",  -- 129
        49440 => X"89",  -- 137
        49441 => X"B1",  -- 177
        49442 => X"AD",  -- 173
        49443 => X"B3",  -- 179
        49444 => X"AB",  -- 171
        49445 => X"96",  -- 150
        49446 => X"9B",  -- 155
        49447 => X"A2",  -- 162
        49448 => X"B9",  -- 185
        49449 => X"97",  -- 151
        49450 => X"62",  -- 98
        49451 => X"3A",  -- 58
        49452 => X"3A",  -- 58
        49453 => X"1E",  -- 30
        49454 => X"28",  -- 40
        49455 => X"31",  -- 49
        49456 => X"34",  -- 52
        49457 => X"37",  -- 55
        49458 => X"35",  -- 53
        49459 => X"2F",  -- 47
        49460 => X"2C",  -- 44
        49461 => X"2E",  -- 46
        49462 => X"31",  -- 49
        49463 => X"32",  -- 50
        49464 => X"32",  -- 50
        49465 => X"2A",  -- 42
        49466 => X"2C",  -- 44
        49467 => X"3D",  -- 61
        49468 => X"4C",  -- 76
        49469 => X"4E",  -- 78
        49470 => X"47",  -- 71
        49471 => X"42",  -- 66
        49472 => X"40",  -- 64
        49473 => X"3C",  -- 60
        49474 => X"3B",  -- 59
        49475 => X"3B",  -- 59
        49476 => X"3A",  -- 58
        49477 => X"37",  -- 55
        49478 => X"36",  -- 54
        49479 => X"38",  -- 56
        49480 => X"36",  -- 54
        49481 => X"30",  -- 48
        49482 => X"2C",  -- 44
        49483 => X"30",  -- 48
        49484 => X"35",  -- 53
        49485 => X"37",  -- 55
        49486 => X"38",  -- 56
        49487 => X"39",  -- 57
        49488 => X"3A",  -- 58
        49489 => X"3B",  -- 59
        49490 => X"37",  -- 55
        49491 => X"35",  -- 53
        49492 => X"39",  -- 57
        49493 => X"41",  -- 65
        49494 => X"45",  -- 69
        49495 => X"45",  -- 69
        49496 => X"47",  -- 71
        49497 => X"44",  -- 68
        49498 => X"48",  -- 72
        49499 => X"48",  -- 72
        49500 => X"41",  -- 65
        49501 => X"41",  -- 65
        49502 => X"48",  -- 72
        49503 => X"4B",  -- 75
        49504 => X"5E",  -- 94
        49505 => X"82",  -- 130
        49506 => X"9B",  -- 155
        49507 => X"9C",  -- 156
        49508 => X"9B",  -- 155
        49509 => X"99",  -- 153
        49510 => X"93",  -- 147
        49511 => X"90",  -- 144
        49512 => X"8B",  -- 139
        49513 => X"8C",  -- 140
        49514 => X"8C",  -- 140
        49515 => X"8D",  -- 141
        49516 => X"93",  -- 147
        49517 => X"9B",  -- 155
        49518 => X"9E",  -- 158
        49519 => X"9F",  -- 159
        49520 => X"A4",  -- 164
        49521 => X"9A",  -- 154
        49522 => X"A3",  -- 163
        49523 => X"AD",  -- 173
        49524 => X"BA",  -- 186
        49525 => X"A6",  -- 166
        49526 => X"A2",  -- 162
        49527 => X"9E",  -- 158
        49528 => X"9B",  -- 155
        49529 => X"9A",  -- 154
        49530 => X"9A",  -- 154
        49531 => X"A1",  -- 161
        49532 => X"9B",  -- 155
        49533 => X"9D",  -- 157
        49534 => X"AB",  -- 171
        49535 => X"9D",  -- 157
        49536 => X"A1",  -- 161
        49537 => X"9F",  -- 159
        49538 => X"A0",  -- 160
        49539 => X"A8",  -- 168
        49540 => X"AC",  -- 172
        49541 => X"A7",  -- 167
        49542 => X"A6",  -- 166
        49543 => X"A8",  -- 168
        49544 => X"B1",  -- 177
        49545 => X"AE",  -- 174
        49546 => X"B2",  -- 178
        49547 => X"BA",  -- 186
        49548 => X"BA",  -- 186
        49549 => X"B5",  -- 181
        49550 => X"B7",  -- 183
        49551 => X"BE",  -- 190
        49552 => X"BA",  -- 186
        49553 => X"B9",  -- 185
        49554 => X"B5",  -- 181
        49555 => X"AF",  -- 175
        49556 => X"B3",  -- 179
        49557 => X"BC",  -- 188
        49558 => X"C1",  -- 193
        49559 => X"BD",  -- 189
        49560 => X"B6",  -- 182
        49561 => X"B5",  -- 181
        49562 => X"B7",  -- 183
        49563 => X"BC",  -- 188
        49564 => X"C0",  -- 192
        49565 => X"C1",  -- 193
        49566 => X"C4",  -- 196
        49567 => X"C7",  -- 199
        49568 => X"C5",  -- 197
        49569 => X"C1",  -- 193
        49570 => X"C1",  -- 193
        49571 => X"C4",  -- 196
        49572 => X"C6",  -- 198
        49573 => X"C4",  -- 196
        49574 => X"C0",  -- 192
        49575 => X"C0",  -- 192
        49576 => X"C1",  -- 193
        49577 => X"A9",  -- 169
        49578 => X"9F",  -- 159
        49579 => X"9F",  -- 159
        49580 => X"95",  -- 149
        49581 => X"82",  -- 130
        49582 => X"6D",  -- 109
        49583 => X"5B",  -- 91
        49584 => X"72",  -- 114
        49585 => X"5F",  -- 95
        49586 => X"44",  -- 68
        49587 => X"3A",  -- 58
        49588 => X"40",  -- 64
        49589 => X"41",  -- 65
        49590 => X"3C",  -- 60
        49591 => X"3D",  -- 61
        49592 => X"44",  -- 68
        49593 => X"51",  -- 81
        49594 => X"5E",  -- 94
        49595 => X"66",  -- 102
        49596 => X"71",  -- 113
        49597 => X"86",  -- 134
        49598 => X"98",  -- 152
        49599 => X"A0",  -- 160
        49600 => X"3A",  -- 58
        49601 => X"3D",  -- 61
        49602 => X"40",  -- 64
        49603 => X"3F",  -- 63
        49604 => X"3C",  -- 60
        49605 => X"3A",  -- 58
        49606 => X"3A",  -- 58
        49607 => X"3B",  -- 59
        49608 => X"42",  -- 66
        49609 => X"43",  -- 67
        49610 => X"45",  -- 69
        49611 => X"45",  -- 69
        49612 => X"44",  -- 68
        49613 => X"44",  -- 68
        49614 => X"47",  -- 71
        49615 => X"4A",  -- 74
        49616 => X"46",  -- 70
        49617 => X"49",  -- 73
        49618 => X"4B",  -- 75
        49619 => X"47",  -- 71
        49620 => X"40",  -- 64
        49621 => X"3F",  -- 63
        49622 => X"44",  -- 68
        49623 => X"4B",  -- 75
        49624 => X"4A",  -- 74
        49625 => X"47",  -- 71
        49626 => X"42",  -- 66
        49627 => X"40",  -- 64
        49628 => X"3F",  -- 63
        49629 => X"3D",  -- 61
        49630 => X"3A",  -- 58
        49631 => X"37",  -- 55
        49632 => X"38",  -- 56
        49633 => X"34",  -- 52
        49634 => X"38",  -- 56
        49635 => X"3D",  -- 61
        49636 => X"40",  -- 64
        49637 => X"45",  -- 69
        49638 => X"44",  -- 68
        49639 => X"3F",  -- 63
        49640 => X"53",  -- 83
        49641 => X"67",  -- 103
        49642 => X"62",  -- 98
        49643 => X"4D",  -- 77
        49644 => X"4A",  -- 74
        49645 => X"5D",  -- 93
        49646 => X"5E",  -- 94
        49647 => X"43",  -- 67
        49648 => X"4C",  -- 76
        49649 => X"47",  -- 71
        49650 => X"44",  -- 68
        49651 => X"22",  -- 34
        49652 => X"24",  -- 36
        49653 => X"1F",  -- 31
        49654 => X"17",  -- 23
        49655 => X"14",  -- 20
        49656 => X"18",  -- 24
        49657 => X"27",  -- 39
        49658 => X"5B",  -- 91
        49659 => X"3F",  -- 63
        49660 => X"50",  -- 80
        49661 => X"72",  -- 114
        49662 => X"67",  -- 103
        49663 => X"55",  -- 85
        49664 => X"52",  -- 82
        49665 => X"4B",  -- 75
        49666 => X"45",  -- 69
        49667 => X"3F",  -- 63
        49668 => X"45",  -- 69
        49669 => X"40",  -- 64
        49670 => X"30",  -- 48
        49671 => X"36",  -- 54
        49672 => X"45",  -- 69
        49673 => X"34",  -- 52
        49674 => X"26",  -- 38
        49675 => X"2D",  -- 45
        49676 => X"40",  -- 64
        49677 => X"45",  -- 69
        49678 => X"40",  -- 64
        49679 => X"41",  -- 65
        49680 => X"50",  -- 80
        49681 => X"5B",  -- 91
        49682 => X"69",  -- 105
        49683 => X"72",  -- 114
        49684 => X"6A",  -- 106
        49685 => X"78",  -- 120
        49686 => X"70",  -- 112
        49687 => X"7D",  -- 125
        49688 => X"87",  -- 135
        49689 => X"85",  -- 133
        49690 => X"81",  -- 129
        49691 => X"89",  -- 137
        49692 => X"95",  -- 149
        49693 => X"90",  -- 144
        49694 => X"85",  -- 133
        49695 => X"84",  -- 132
        49696 => X"79",  -- 121
        49697 => X"88",  -- 136
        49698 => X"84",  -- 132
        49699 => X"7A",  -- 122
        49700 => X"82",  -- 130
        49701 => X"7C",  -- 124
        49702 => X"7B",  -- 123
        49703 => X"87",  -- 135
        49704 => X"81",  -- 129
        49705 => X"73",  -- 115
        49706 => X"6F",  -- 111
        49707 => X"76",  -- 118
        49708 => X"6D",  -- 109
        49709 => X"58",  -- 88
        49710 => X"52",  -- 82
        49711 => X"52",  -- 82
        49712 => X"57",  -- 87
        49713 => X"5C",  -- 92
        49714 => X"64",  -- 100
        49715 => X"6F",  -- 111
        49716 => X"78",  -- 120
        49717 => X"7B",  -- 123
        49718 => X"7B",  -- 123
        49719 => X"79",  -- 121
        49720 => X"6E",  -- 110
        49721 => X"6B",  -- 107
        49722 => X"81",  -- 129
        49723 => X"8D",  -- 141
        49724 => X"82",  -- 130
        49725 => X"90",  -- 144
        49726 => X"9E",  -- 158
        49727 => X"91",  -- 145
        49728 => X"75",  -- 117
        49729 => X"8B",  -- 139
        49730 => X"D7",  -- 215
        49731 => X"83",  -- 131
        49732 => X"9A",  -- 154
        49733 => X"C4",  -- 196
        49734 => X"96",  -- 150
        49735 => X"86",  -- 134
        49736 => X"6B",  -- 107
        49737 => X"5D",  -- 93
        49738 => X"6B",  -- 107
        49739 => X"43",  -- 67
        49740 => X"0A",  -- 10
        49741 => X"0B",  -- 11
        49742 => X"0D",  -- 13
        49743 => X"05",  -- 5
        49744 => X"18",  -- 24
        49745 => X"29",  -- 41
        49746 => X"3B",  -- 59
        49747 => X"52",  -- 82
        49748 => X"5F",  -- 95
        49749 => X"74",  -- 116
        49750 => X"6A",  -- 106
        49751 => X"62",  -- 98
        49752 => X"67",  -- 103
        49753 => X"7C",  -- 124
        49754 => X"91",  -- 145
        49755 => X"A9",  -- 169
        49756 => X"8D",  -- 141
        49757 => X"A1",  -- 161
        49758 => X"84",  -- 132
        49759 => X"81",  -- 129
        49760 => X"8C",  -- 140
        49761 => X"B1",  -- 177
        49762 => X"B1",  -- 177
        49763 => X"B9",  -- 185
        49764 => X"AC",  -- 172
        49765 => X"9C",  -- 156
        49766 => X"93",  -- 147
        49767 => X"91",  -- 145
        49768 => X"AD",  -- 173
        49769 => X"A5",  -- 165
        49770 => X"6D",  -- 109
        49771 => X"27",  -- 39
        49772 => X"2D",  -- 45
        49773 => X"2A",  -- 42
        49774 => X"37",  -- 55
        49775 => X"2D",  -- 45
        49776 => X"35",  -- 53
        49777 => X"38",  -- 56
        49778 => X"35",  -- 53
        49779 => X"2F",  -- 47
        49780 => X"2C",  -- 44
        49781 => X"2D",  -- 45
        49782 => X"30",  -- 48
        49783 => X"30",  -- 48
        49784 => X"2E",  -- 46
        49785 => X"29",  -- 41
        49786 => X"2C",  -- 44
        49787 => X"3C",  -- 60
        49788 => X"4B",  -- 75
        49789 => X"4F",  -- 79
        49790 => X"49",  -- 73
        49791 => X"43",  -- 67
        49792 => X"41",  -- 65
        49793 => X"3E",  -- 62
        49794 => X"3C",  -- 60
        49795 => X"3B",  -- 59
        49796 => X"3B",  -- 59
        49797 => X"39",  -- 57
        49798 => X"38",  -- 56
        49799 => X"37",  -- 55
        49800 => X"36",  -- 54
        49801 => X"2F",  -- 47
        49802 => X"2B",  -- 43
        49803 => X"2F",  -- 47
        49804 => X"35",  -- 53
        49805 => X"37",  -- 55
        49806 => X"38",  -- 56
        49807 => X"38",  -- 56
        49808 => X"3C",  -- 60
        49809 => X"3E",  -- 62
        49810 => X"3C",  -- 60
        49811 => X"37",  -- 55
        49812 => X"37",  -- 55
        49813 => X"3F",  -- 63
        49814 => X"45",  -- 69
        49815 => X"48",  -- 72
        49816 => X"47",  -- 71
        49817 => X"43",  -- 67
        49818 => X"48",  -- 72
        49819 => X"49",  -- 73
        49820 => X"3E",  -- 62
        49821 => X"3F",  -- 63
        49822 => X"52",  -- 82
        49823 => X"63",  -- 99
        49824 => X"8A",  -- 138
        49825 => X"A6",  -- 166
        49826 => X"A9",  -- 169
        49827 => X"9E",  -- 158
        49828 => X"9C",  -- 156
        49829 => X"99",  -- 153
        49830 => X"93",  -- 147
        49831 => X"98",  -- 152
        49832 => X"93",  -- 147
        49833 => X"93",  -- 147
        49834 => X"90",  -- 144
        49835 => X"91",  -- 145
        49836 => X"9A",  -- 154
        49837 => X"A5",  -- 165
        49838 => X"A7",  -- 167
        49839 => X"A2",  -- 162
        49840 => X"B1",  -- 177
        49841 => X"A8",  -- 168
        49842 => X"AD",  -- 173
        49843 => X"A8",  -- 168
        49844 => X"AE",  -- 174
        49845 => X"A7",  -- 167
        49846 => X"B1",  -- 177
        49847 => X"AB",  -- 171
        49848 => X"AB",  -- 171
        49849 => X"A4",  -- 164
        49850 => X"A5",  -- 165
        49851 => X"A9",  -- 169
        49852 => X"99",  -- 153
        49853 => X"99",  -- 153
        49854 => X"A8",  -- 168
        49855 => X"94",  -- 148
        49856 => X"A4",  -- 164
        49857 => X"A0",  -- 160
        49858 => X"A4",  -- 164
        49859 => X"B0",  -- 176
        49860 => X"B2",  -- 178
        49861 => X"AD",  -- 173
        49862 => X"AB",  -- 171
        49863 => X"AF",  -- 175
        49864 => X"AE",  -- 174
        49865 => X"A8",  -- 168
        49866 => X"AE",  -- 174
        49867 => X"BA",  -- 186
        49868 => X"BD",  -- 189
        49869 => X"B3",  -- 179
        49870 => X"B3",  -- 179
        49871 => X"BC",  -- 188
        49872 => X"B9",  -- 185
        49873 => X"B5",  -- 181
        49874 => X"AD",  -- 173
        49875 => X"AC",  -- 172
        49876 => X"B6",  -- 182
        49877 => X"C0",  -- 192
        49878 => X"C1",  -- 193
        49879 => X"BA",  -- 186
        49880 => X"B9",  -- 185
        49881 => X"B6",  -- 182
        49882 => X"B5",  -- 181
        49883 => X"B9",  -- 185
        49884 => X"C0",  -- 192
        49885 => X"C4",  -- 196
        49886 => X"C6",  -- 198
        49887 => X"C6",  -- 198
        49888 => X"C6",  -- 198
        49889 => X"C1",  -- 193
        49890 => X"BF",  -- 191
        49891 => X"C2",  -- 194
        49892 => X"C4",  -- 196
        49893 => X"C2",  -- 194
        49894 => X"BF",  -- 191
        49895 => X"BF",  -- 191
        49896 => X"B6",  -- 182
        49897 => X"B4",  -- 180
        49898 => X"A6",  -- 166
        49899 => X"8D",  -- 141
        49900 => X"88",  -- 136
        49901 => X"93",  -- 147
        49902 => X"7E",  -- 126
        49903 => X"4F",  -- 79
        49904 => X"55",  -- 85
        49905 => X"55",  -- 85
        49906 => X"3F",  -- 63
        49907 => X"2C",  -- 44
        49908 => X"31",  -- 49
        49909 => X"36",  -- 54
        49910 => X"3C",  -- 60
        49911 => X"4D",  -- 77
        49912 => X"42",  -- 66
        49913 => X"50",  -- 80
        49914 => X"63",  -- 99
        49915 => X"71",  -- 113
        49916 => X"7D",  -- 125
        49917 => X"8B",  -- 139
        49918 => X"95",  -- 149
        49919 => X"9B",  -- 155
        49920 => X"39",  -- 57
        49921 => X"3B",  -- 59
        49922 => X"3C",  -- 60
        49923 => X"3A",  -- 58
        49924 => X"37",  -- 55
        49925 => X"37",  -- 55
        49926 => X"3A",  -- 58
        49927 => X"3E",  -- 62
        49928 => X"3B",  -- 59
        49929 => X"3C",  -- 60
        49930 => X"3D",  -- 61
        49931 => X"3D",  -- 61
        49932 => X"3E",  -- 62
        49933 => X"3F",  -- 63
        49934 => X"41",  -- 65
        49935 => X"44",  -- 68
        49936 => X"3E",  -- 62
        49937 => X"3F",  -- 63
        49938 => X"3F",  -- 63
        49939 => X"3D",  -- 61
        49940 => X"3D",  -- 61
        49941 => X"3C",  -- 60
        49942 => X"3E",  -- 62
        49943 => X"40",  -- 64
        49944 => X"41",  -- 65
        49945 => X"3E",  -- 62
        49946 => X"3C",  -- 60
        49947 => X"3C",  -- 60
        49948 => X"3C",  -- 60
        49949 => X"3A",  -- 58
        49950 => X"36",  -- 54
        49951 => X"32",  -- 50
        49952 => X"31",  -- 49
        49953 => X"31",  -- 49
        49954 => X"31",  -- 49
        49955 => X"35",  -- 53
        49956 => X"3C",  -- 60
        49957 => X"3D",  -- 61
        49958 => X"37",  -- 55
        49959 => X"35",  -- 53
        49960 => X"58",  -- 88
        49961 => X"61",  -- 97
        49962 => X"5C",  -- 92
        49963 => X"49",  -- 73
        49964 => X"52",  -- 82
        49965 => X"65",  -- 101
        49966 => X"55",  -- 85
        49967 => X"39",  -- 57
        49968 => X"54",  -- 84
        49969 => X"55",  -- 85
        49970 => X"53",  -- 83
        49971 => X"31",  -- 49
        49972 => X"31",  -- 49
        49973 => X"29",  -- 41
        49974 => X"1D",  -- 29
        49975 => X"16",  -- 22
        49976 => X"1A",  -- 26
        49977 => X"22",  -- 34
        49978 => X"4C",  -- 76
        49979 => X"5B",  -- 91
        49980 => X"6F",  -- 111
        49981 => X"6D",  -- 109
        49982 => X"68",  -- 104
        49983 => X"57",  -- 87
        49984 => X"4A",  -- 74
        49985 => X"45",  -- 69
        49986 => X"49",  -- 73
        49987 => X"44",  -- 68
        49988 => X"44",  -- 68
        49989 => X"43",  -- 67
        49990 => X"36",  -- 54
        49991 => X"3B",  -- 59
        49992 => X"3F",  -- 63
        49993 => X"31",  -- 49
        49994 => X"20",  -- 32
        49995 => X"2B",  -- 43
        49996 => X"48",  -- 72
        49997 => X"4F",  -- 79
        49998 => X"47",  -- 71
        49999 => X"48",  -- 72
        50000 => X"52",  -- 82
        50001 => X"5A",  -- 90
        50002 => X"69",  -- 105
        50003 => X"74",  -- 116
        50004 => X"6F",  -- 111
        50005 => X"7B",  -- 123
        50006 => X"73",  -- 115
        50007 => X"80",  -- 128
        50008 => X"85",  -- 133
        50009 => X"82",  -- 130
        50010 => X"7C",  -- 124
        50011 => X"80",  -- 128
        50012 => X"8B",  -- 139
        50013 => X"8A",  -- 138
        50014 => X"80",  -- 128
        50015 => X"7E",  -- 126
        50016 => X"81",  -- 129
        50017 => X"8D",  -- 141
        50018 => X"95",  -- 149
        50019 => X"75",  -- 117
        50020 => X"83",  -- 131
        50021 => X"7B",  -- 123
        50022 => X"8C",  -- 140
        50023 => X"8F",  -- 143
        50024 => X"7F",  -- 127
        50025 => X"71",  -- 113
        50026 => X"78",  -- 120
        50027 => X"7B",  -- 123
        50028 => X"65",  -- 101
        50029 => X"51",  -- 81
        50030 => X"48",  -- 72
        50031 => X"49",  -- 73
        50032 => X"65",  -- 101
        50033 => X"74",  -- 116
        50034 => X"7E",  -- 126
        50035 => X"79",  -- 121
        50036 => X"78",  -- 120
        50037 => X"83",  -- 131
        50038 => X"85",  -- 133
        50039 => X"7D",  -- 125
        50040 => X"76",  -- 118
        50041 => X"75",  -- 117
        50042 => X"7A",  -- 122
        50043 => X"82",  -- 130
        50044 => X"88",  -- 136
        50045 => X"99",  -- 153
        50046 => X"B0",  -- 176
        50047 => X"BF",  -- 191
        50048 => X"9F",  -- 159
        50049 => X"6E",  -- 110
        50050 => X"CA",  -- 202
        50051 => X"A8",  -- 168
        50052 => X"9F",  -- 159
        50053 => X"A7",  -- 167
        50054 => X"6E",  -- 110
        50055 => X"5D",  -- 93
        50056 => X"4A",  -- 74
        50057 => X"33",  -- 51
        50058 => X"4A",  -- 74
        50059 => X"3C",  -- 60
        50060 => X"15",  -- 21
        50061 => X"12",  -- 18
        50062 => X"14",  -- 20
        50063 => X"14",  -- 20
        50064 => X"28",  -- 40
        50065 => X"3E",  -- 62
        50066 => X"48",  -- 72
        50067 => X"64",  -- 100
        50068 => X"67",  -- 103
        50069 => X"77",  -- 119
        50070 => X"6F",  -- 111
        50071 => X"6A",  -- 106
        50072 => X"6F",  -- 111
        50073 => X"77",  -- 119
        50074 => X"8E",  -- 142
        50075 => X"AA",  -- 170
        50076 => X"8D",  -- 141
        50077 => X"9A",  -- 154
        50078 => X"88",  -- 136
        50079 => X"7E",  -- 126
        50080 => X"92",  -- 146
        50081 => X"B1",  -- 177
        50082 => X"B0",  -- 176
        50083 => X"B9",  -- 185
        50084 => X"A7",  -- 167
        50085 => X"A3",  -- 163
        50086 => X"93",  -- 147
        50087 => X"89",  -- 137
        50088 => X"9A",  -- 154
        50089 => X"9D",  -- 157
        50090 => X"61",  -- 97
        50091 => X"20",  -- 32
        50092 => X"2B",  -- 43
        50093 => X"36",  -- 54
        50094 => X"41",  -- 65
        50095 => X"37",  -- 55
        50096 => X"36",  -- 54
        50097 => X"37",  -- 55
        50098 => X"34",  -- 52
        50099 => X"2E",  -- 46
        50100 => X"2B",  -- 43
        50101 => X"2F",  -- 47
        50102 => X"31",  -- 49
        50103 => X"30",  -- 48
        50104 => X"2D",  -- 45
        50105 => X"28",  -- 40
        50106 => X"2B",  -- 43
        50107 => X"39",  -- 57
        50108 => X"48",  -- 72
        50109 => X"4D",  -- 77
        50110 => X"4A",  -- 74
        50111 => X"44",  -- 68
        50112 => X"42",  -- 66
        50113 => X"40",  -- 64
        50114 => X"3E",  -- 62
        50115 => X"3C",  -- 60
        50116 => X"3C",  -- 60
        50117 => X"3B",  -- 59
        50118 => X"39",  -- 57
        50119 => X"36",  -- 54
        50120 => X"35",  -- 53
        50121 => X"2F",  -- 47
        50122 => X"2D",  -- 45
        50123 => X"31",  -- 49
        50124 => X"36",  -- 54
        50125 => X"37",  -- 55
        50126 => X"37",  -- 55
        50127 => X"38",  -- 56
        50128 => X"3A",  -- 58
        50129 => X"40",  -- 64
        50130 => X"41",  -- 65
        50131 => X"3D",  -- 61
        50132 => X"3A",  -- 58
        50133 => X"3F",  -- 63
        50134 => X"4A",  -- 74
        50135 => X"50",  -- 80
        50136 => X"48",  -- 72
        50137 => X"47",  -- 71
        50138 => X"4C",  -- 76
        50139 => X"4B",  -- 75
        50140 => X"41",  -- 65
        50141 => X"4B",  -- 75
        50142 => X"6D",  -- 109
        50143 => X"89",  -- 137
        50144 => X"9E",  -- 158
        50145 => X"A3",  -- 163
        50146 => X"99",  -- 153
        50147 => X"96",  -- 150
        50148 => X"9E",  -- 158
        50149 => X"9B",  -- 155
        50150 => X"98",  -- 152
        50151 => X"A6",  -- 166
        50152 => X"9F",  -- 159
        50153 => X"97",  -- 151
        50154 => X"90",  -- 144
        50155 => X"93",  -- 147
        50156 => X"A1",  -- 161
        50157 => X"AC",  -- 172
        50158 => X"AB",  -- 171
        50159 => X"A4",  -- 164
        50160 => X"B6",  -- 182
        50161 => X"B4",  -- 180
        50162 => X"BC",  -- 188
        50163 => X"A9",  -- 169
        50164 => X"A4",  -- 164
        50165 => X"A7",  -- 167
        50166 => X"B7",  -- 183
        50167 => X"AE",  -- 174
        50168 => X"A6",  -- 166
        50169 => X"A1",  -- 161
        50170 => X"A2",  -- 162
        50171 => X"A8",  -- 168
        50172 => X"99",  -- 153
        50173 => X"9A",  -- 154
        50174 => X"A9",  -- 169
        50175 => X"93",  -- 147
        50176 => X"A5",  -- 165
        50177 => X"A3",  -- 163
        50178 => X"A9",  -- 169
        50179 => X"B3",  -- 179
        50180 => X"B7",  -- 183
        50181 => X"B3",  -- 179
        50182 => X"B1",  -- 177
        50183 => X"B3",  -- 179
        50184 => X"B1",  -- 177
        50185 => X"A6",  -- 166
        50186 => X"A9",  -- 169
        50187 => X"B8",  -- 184
        50188 => X"BE",  -- 190
        50189 => X"B3",  -- 179
        50190 => X"B0",  -- 176
        50191 => X"B6",  -- 182
        50192 => X"BA",  -- 186
        50193 => X"B1",  -- 177
        50194 => X"A9",  -- 169
        50195 => X"AC",  -- 172
        50196 => X"BB",  -- 187
        50197 => X"C5",  -- 197
        50198 => X"C3",  -- 195
        50199 => X"BB",  -- 187
        50200 => X"BB",  -- 187
        50201 => X"B9",  -- 185
        50202 => X"B8",  -- 184
        50203 => X"BA",  -- 186
        50204 => X"C0",  -- 192
        50205 => X"C5",  -- 197
        50206 => X"C6",  -- 198
        50207 => X"C5",  -- 197
        50208 => X"C7",  -- 199
        50209 => X"C2",  -- 194
        50210 => X"BF",  -- 191
        50211 => X"C1",  -- 193
        50212 => X"C3",  -- 195
        50213 => X"C0",  -- 192
        50214 => X"BE",  -- 190
        50215 => X"BE",  -- 190
        50216 => X"BD",  -- 189
        50217 => X"AE",  -- 174
        50218 => X"9F",  -- 159
        50219 => X"91",  -- 145
        50220 => X"87",  -- 135
        50221 => X"86",  -- 134
        50222 => X"7E",  -- 126
        50223 => X"6A",  -- 106
        50224 => X"49",  -- 73
        50225 => X"50",  -- 80
        50226 => X"40",  -- 64
        50227 => X"29",  -- 41
        50228 => X"2A",  -- 42
        50229 => X"30",  -- 48
        50230 => X"3B",  -- 59
        50231 => X"4F",  -- 79
        50232 => X"49",  -- 73
        50233 => X"4D",  -- 77
        50234 => X"61",  -- 97
        50235 => X"7D",  -- 125
        50236 => X"8F",  -- 143
        50237 => X"94",  -- 148
        50238 => X"99",  -- 153
        50239 => X"A0",  -- 160
        50240 => X"3F",  -- 63
        50241 => X"3E",  -- 62
        50242 => X"3D",  -- 61
        50243 => X"3C",  -- 60
        50244 => X"3C",  -- 60
        50245 => X"3E",  -- 62
        50246 => X"42",  -- 66
        50247 => X"45",  -- 69
        50248 => X"41",  -- 65
        50249 => X"3F",  -- 63
        50250 => X"3D",  -- 61
        50251 => X"3E",  -- 62
        50252 => X"41",  -- 65
        50253 => X"44",  -- 68
        50254 => X"46",  -- 70
        50255 => X"47",  -- 71
        50256 => X"42",  -- 66
        50257 => X"41",  -- 65
        50258 => X"3F",  -- 63
        50259 => X"40",  -- 64
        50260 => X"43",  -- 67
        50261 => X"43",  -- 67
        50262 => X"40",  -- 64
        50263 => X"3E",  -- 62
        50264 => X"3A",  -- 58
        50265 => X"39",  -- 57
        50266 => X"3A",  -- 58
        50267 => X"3B",  -- 59
        50268 => X"3C",  -- 60
        50269 => X"39",  -- 57
        50270 => X"34",  -- 52
        50271 => X"30",  -- 48
        50272 => X"2D",  -- 45
        50273 => X"31",  -- 49
        50274 => X"2F",  -- 47
        50275 => X"34",  -- 52
        50276 => X"3D",  -- 61
        50277 => X"3B",  -- 59
        50278 => X"34",  -- 52
        50279 => X"38",  -- 56
        50280 => X"5D",  -- 93
        50281 => X"5B",  -- 91
        50282 => X"54",  -- 84
        50283 => X"45",  -- 69
        50284 => X"57",  -- 87
        50285 => X"67",  -- 103
        50286 => X"4B",  -- 75
        50287 => X"34",  -- 52
        50288 => X"53",  -- 83
        50289 => X"56",  -- 86
        50290 => X"5A",  -- 90
        50291 => X"3C",  -- 60
        50292 => X"3D",  -- 61
        50293 => X"33",  -- 51
        50294 => X"28",  -- 40
        50295 => X"24",  -- 36
        50296 => X"22",  -- 34
        50297 => X"24",  -- 36
        50298 => X"3C",  -- 60
        50299 => X"71",  -- 113
        50300 => X"85",  -- 133
        50301 => X"6D",  -- 109
        50302 => X"6C",  -- 108
        50303 => X"5E",  -- 94
        50304 => X"4D",  -- 77
        50305 => X"49",  -- 73
        50306 => X"50",  -- 80
        50307 => X"4A",  -- 74
        50308 => X"45",  -- 69
        50309 => X"44",  -- 68
        50310 => X"3B",  -- 59
        50311 => X"3D",  -- 61
        50312 => X"3D",  -- 61
        50313 => X"2C",  -- 44
        50314 => X"15",  -- 21
        50315 => X"20",  -- 32
        50316 => X"47",  -- 71
        50317 => X"52",  -- 82
        50318 => X"47",  -- 71
        50319 => X"48",  -- 72
        50320 => X"4C",  -- 76
        50321 => X"53",  -- 83
        50322 => X"63",  -- 99
        50323 => X"72",  -- 114
        50324 => X"6E",  -- 110
        50325 => X"78",  -- 120
        50326 => X"6B",  -- 107
        50327 => X"75",  -- 117
        50328 => X"80",  -- 128
        50329 => X"87",  -- 135
        50330 => X"86",  -- 134
        50331 => X"81",  -- 129
        50332 => X"82",  -- 130
        50333 => X"7F",  -- 127
        50334 => X"7C",  -- 124
        50335 => X"80",  -- 128
        50336 => X"8E",  -- 142
        50337 => X"8D",  -- 141
        50338 => X"9C",  -- 156
        50339 => X"7B",  -- 123
        50340 => X"84",  -- 132
        50341 => X"78",  -- 120
        50342 => X"8F",  -- 143
        50343 => X"87",  -- 135
        50344 => X"87",  -- 135
        50345 => X"7E",  -- 126
        50346 => X"87",  -- 135
        50347 => X"79",  -- 121
        50348 => X"66",  -- 102
        50349 => X"66",  -- 102
        50350 => X"4F",  -- 79
        50351 => X"33",  -- 51
        50352 => X"56",  -- 86
        50353 => X"73",  -- 115
        50354 => X"81",  -- 129
        50355 => X"78",  -- 120
        50356 => X"75",  -- 117
        50357 => X"83",  -- 131
        50358 => X"8A",  -- 138
        50359 => X"85",  -- 133
        50360 => X"83",  -- 131
        50361 => X"8B",  -- 139
        50362 => X"84",  -- 132
        50363 => X"7D",  -- 125
        50364 => X"8C",  -- 140
        50365 => X"A3",  -- 163
        50366 => X"B0",  -- 176
        50367 => X"B6",  -- 182
        50368 => X"A9",  -- 169
        50369 => X"74",  -- 116
        50370 => X"BC",  -- 188
        50371 => X"B4",  -- 180
        50372 => X"88",  -- 136
        50373 => X"71",  -- 113
        50374 => X"43",  -- 67
        50375 => X"37",  -- 55
        50376 => X"31",  -- 49
        50377 => X"18",  -- 24
        50378 => X"25",  -- 37
        50379 => X"2B",  -- 43
        50380 => X"17",  -- 23
        50381 => X"17",  -- 23
        50382 => X"1F",  -- 31
        50383 => X"23",  -- 35
        50384 => X"35",  -- 53
        50385 => X"4E",  -- 78
        50386 => X"4E",  -- 78
        50387 => X"6B",  -- 107
        50388 => X"66",  -- 102
        50389 => X"76",  -- 118
        50390 => X"75",  -- 117
        50391 => X"75",  -- 117
        50392 => X"71",  -- 113
        50393 => X"6E",  -- 110
        50394 => X"86",  -- 134
        50395 => X"A4",  -- 164
        50396 => X"90",  -- 144
        50397 => X"8D",  -- 141
        50398 => X"86",  -- 134
        50399 => X"79",  -- 121
        50400 => X"95",  -- 149
        50401 => X"AD",  -- 173
        50402 => X"AB",  -- 171
        50403 => X"B3",  -- 179
        50404 => X"9D",  -- 157
        50405 => X"A6",  -- 166
        50406 => X"90",  -- 144
        50407 => X"83",  -- 131
        50408 => X"90",  -- 144
        50409 => X"8A",  -- 138
        50410 => X"45",  -- 69
        50411 => X"20",  -- 32
        50412 => X"2C",  -- 44
        50413 => X"33",  -- 51
        50414 => X"33",  -- 51
        50415 => X"39",  -- 57
        50416 => X"38",  -- 56
        50417 => X"37",  -- 55
        50418 => X"34",  -- 52
        50419 => X"2E",  -- 46
        50420 => X"2D",  -- 45
        50421 => X"2F",  -- 47
        50422 => X"31",  -- 49
        50423 => X"30",  -- 48
        50424 => X"2E",  -- 46
        50425 => X"2B",  -- 43
        50426 => X"2C",  -- 44
        50427 => X"37",  -- 55
        50428 => X"45",  -- 69
        50429 => X"4C",  -- 76
        50430 => X"4B",  -- 75
        50431 => X"45",  -- 69
        50432 => X"42",  -- 66
        50433 => X"41",  -- 65
        50434 => X"3F",  -- 63
        50435 => X"3D",  -- 61
        50436 => X"3D",  -- 61
        50437 => X"3E",  -- 62
        50438 => X"3A",  -- 58
        50439 => X"35",  -- 53
        50440 => X"32",  -- 50
        50441 => X"30",  -- 48
        50442 => X"30",  -- 48
        50443 => X"35",  -- 53
        50444 => X"38",  -- 56
        50445 => X"37",  -- 55
        50446 => X"37",  -- 55
        50447 => X"39",  -- 57
        50448 => X"40",  -- 64
        50449 => X"45",  -- 69
        50450 => X"45",  -- 69
        50451 => X"3E",  -- 62
        50452 => X"38",  -- 56
        50453 => X"3C",  -- 60
        50454 => X"44",  -- 68
        50455 => X"4A",  -- 74
        50456 => X"46",  -- 70
        50457 => X"46",  -- 70
        50458 => X"4C",  -- 76
        50459 => X"4B",  -- 75
        50460 => X"46",  -- 70
        50461 => X"59",  -- 89
        50462 => X"83",  -- 131
        50463 => X"A0",  -- 160
        50464 => X"91",  -- 145
        50465 => X"86",  -- 134
        50466 => X"81",  -- 129
        50467 => X"8C",  -- 140
        50468 => X"9C",  -- 156
        50469 => X"9B",  -- 155
        50470 => X"9E",  -- 158
        50471 => X"AC",  -- 172
        50472 => X"A9",  -- 169
        50473 => X"9B",  -- 155
        50474 => X"91",  -- 145
        50475 => X"96",  -- 150
        50476 => X"A3",  -- 163
        50477 => X"A8",  -- 168
        50478 => X"A6",  -- 166
        50479 => X"A2",  -- 162
        50480 => X"AE",  -- 174
        50481 => X"AF",  -- 175
        50482 => X"C2",  -- 194
        50483 => X"B1",  -- 177
        50484 => X"A7",  -- 167
        50485 => X"A7",  -- 167
        50486 => X"B8",  -- 184
        50487 => X"A7",  -- 167
        50488 => X"9E",  -- 158
        50489 => X"9E",  -- 158
        50490 => X"A0",  -- 160
        50491 => X"A7",  -- 167
        50492 => X"9F",  -- 159
        50493 => X"A1",  -- 161
        50494 => X"AE",  -- 174
        50495 => X"A0",  -- 160
        50496 => X"A2",  -- 162
        50497 => X"A4",  -- 164
        50498 => X"AA",  -- 170
        50499 => X"AF",  -- 175
        50500 => X"B5",  -- 181
        50501 => X"B7",  -- 183
        50502 => X"B6",  -- 182
        50503 => X"B4",  -- 180
        50504 => X"B7",  -- 183
        50505 => X"AB",  -- 171
        50506 => X"AA",  -- 170
        50507 => X"B7",  -- 183
        50508 => X"BC",  -- 188
        50509 => X"B3",  -- 179
        50510 => X"AE",  -- 174
        50511 => X"B1",  -- 177
        50512 => X"BA",  -- 186
        50513 => X"B2",  -- 178
        50514 => X"AC",  -- 172
        50515 => X"AF",  -- 175
        50516 => X"BB",  -- 187
        50517 => X"C3",  -- 195
        50518 => X"C0",  -- 192
        50519 => X"BA",  -- 186
        50520 => X"B9",  -- 185
        50521 => X"B9",  -- 185
        50522 => X"BB",  -- 187
        50523 => X"BB",  -- 187
        50524 => X"BF",  -- 191
        50525 => X"C4",  -- 196
        50526 => X"C6",  -- 198
        50527 => X"C4",  -- 196
        50528 => X"C8",  -- 200
        50529 => X"C2",  -- 194
        50530 => X"BF",  -- 191
        50531 => X"C1",  -- 193
        50532 => X"C1",  -- 193
        50533 => X"BE",  -- 190
        50534 => X"BB",  -- 187
        50535 => X"BA",  -- 186
        50536 => X"BE",  -- 190
        50537 => X"AC",  -- 172
        50538 => X"9F",  -- 159
        50539 => X"92",  -- 146
        50540 => X"81",  -- 129
        50541 => X"79",  -- 121
        50542 => X"7B",  -- 123
        50543 => X"78",  -- 120
        50544 => X"52",  -- 82
        50545 => X"4E",  -- 78
        50546 => X"3C",  -- 60
        50547 => X"2C",  -- 44
        50548 => X"2D",  -- 45
        50549 => X"34",  -- 52
        50550 => X"3E",  -- 62
        50551 => X"4A",  -- 74
        50552 => X"54",  -- 84
        50553 => X"4F",  -- 79
        50554 => X"5D",  -- 93
        50555 => X"7A",  -- 122
        50556 => X"92",  -- 146
        50557 => X"99",  -- 153
        50558 => X"A0",  -- 160
        50559 => X"AB",  -- 171
        50560 => X"43",  -- 67
        50561 => X"42",  -- 66
        50562 => X"41",  -- 65
        50563 => X"42",  -- 66
        50564 => X"45",  -- 69
        50565 => X"47",  -- 71
        50566 => X"49",  -- 73
        50567 => X"4A",  -- 74
        50568 => X"4A",  -- 74
        50569 => X"45",  -- 69
        50570 => X"41",  -- 65
        50571 => X"42",  -- 66
        50572 => X"48",  -- 72
        50573 => X"4D",  -- 77
        50574 => X"4F",  -- 79
        50575 => X"4E",  -- 78
        50576 => X"48",  -- 72
        50577 => X"46",  -- 70
        50578 => X"45",  -- 69
        50579 => X"45",  -- 69
        50580 => X"47",  -- 71
        50581 => X"46",  -- 70
        50582 => X"43",  -- 67
        50583 => X"40",  -- 64
        50584 => X"3B",  -- 59
        50585 => X"3A",  -- 58
        50586 => X"3A",  -- 58
        50587 => X"3B",  -- 59
        50588 => X"3C",  -- 60
        50589 => X"3B",  -- 59
        50590 => X"36",  -- 54
        50591 => X"32",  -- 50
        50592 => X"2D",  -- 45
        50593 => X"32",  -- 50
        50594 => X"2D",  -- 45
        50595 => X"2F",  -- 47
        50596 => X"39",  -- 57
        50597 => X"36",  -- 54
        50598 => X"32",  -- 50
        50599 => X"3E",  -- 62
        50600 => X"55",  -- 85
        50601 => X"4E",  -- 78
        50602 => X"46",  -- 70
        50603 => X"3D",  -- 61
        50604 => X"56",  -- 86
        50605 => X"63",  -- 99
        50606 => X"44",  -- 68
        50607 => X"38",  -- 56
        50608 => X"4E",  -- 78
        50609 => X"52",  -- 82
        50610 => X"5D",  -- 93
        50611 => X"46",  -- 70
        50612 => X"48",  -- 72
        50613 => X"3C",  -- 60
        50614 => X"35",  -- 53
        50615 => X"37",  -- 55
        50616 => X"2F",  -- 47
        50617 => X"2A",  -- 42
        50618 => X"36",  -- 54
        50619 => X"70",  -- 112
        50620 => X"7F",  -- 127
        50621 => X"71",  -- 113
        50622 => X"66",  -- 102
        50623 => X"5A",  -- 90
        50624 => X"53",  -- 83
        50625 => X"4A",  -- 74
        50626 => X"51",  -- 81
        50627 => X"4D",  -- 77
        50628 => X"48",  -- 72
        50629 => X"4A",  -- 74
        50630 => X"41",  -- 65
        50631 => X"3D",  -- 61
        50632 => X"38",  -- 56
        50633 => X"32",  -- 50
        50634 => X"1F",  -- 31
        50635 => X"25",  -- 37
        50636 => X"47",  -- 71
        50637 => X"4B",  -- 75
        50638 => X"43",  -- 67
        50639 => X"4D",  -- 77
        50640 => X"50",  -- 80
        50641 => X"52",  -- 82
        50642 => X"5C",  -- 92
        50643 => X"6C",  -- 108
        50644 => X"6C",  -- 108
        50645 => X"79",  -- 121
        50646 => X"6F",  -- 111
        50647 => X"7A",  -- 122
        50648 => X"7D",  -- 125
        50649 => X"89",  -- 137
        50650 => X"8A",  -- 138
        50651 => X"84",  -- 132
        50652 => X"83",  -- 131
        50653 => X"81",  -- 129
        50654 => X"7D",  -- 125
        50655 => X"80",  -- 128
        50656 => X"8C",  -- 140
        50657 => X"79",  -- 121
        50658 => X"88",  -- 136
        50659 => X"85",  -- 133
        50660 => X"84",  -- 132
        50661 => X"79",  -- 121
        50662 => X"87",  -- 135
        50663 => X"7A",  -- 122
        50664 => X"82",  -- 130
        50665 => X"77",  -- 119
        50666 => X"83",  -- 131
        50667 => X"74",  -- 116
        50668 => X"64",  -- 100
        50669 => X"6B",  -- 107
        50670 => X"49",  -- 73
        50671 => X"1F",  -- 31
        50672 => X"44",  -- 68
        50673 => X"5F",  -- 95
        50674 => X"74",  -- 116
        50675 => X"75",  -- 117
        50676 => X"73",  -- 115
        50677 => X"7D",  -- 125
        50678 => X"88",  -- 136
        50679 => X"8B",  -- 139
        50680 => X"86",  -- 134
        50681 => X"91",  -- 145
        50682 => X"93",  -- 147
        50683 => X"8C",  -- 140
        50684 => X"90",  -- 144
        50685 => X"A8",  -- 168
        50686 => X"B5",  -- 181
        50687 => X"AF",  -- 175
        50688 => X"B7",  -- 183
        50689 => X"A9",  -- 169
        50690 => X"BA",  -- 186
        50691 => X"B3",  -- 179
        50692 => X"75",  -- 117
        50693 => X"47",  -- 71
        50694 => X"31",  -- 49
        50695 => X"3D",  -- 61
        50696 => X"24",  -- 36
        50697 => X"1D",  -- 29
        50698 => X"1B",  -- 27
        50699 => X"26",  -- 38
        50700 => X"24",  -- 36
        50701 => X"23",  -- 35
        50702 => X"30",  -- 48
        50703 => X"30",  -- 48
        50704 => X"3C",  -- 60
        50705 => X"58",  -- 88
        50706 => X"55",  -- 85
        50707 => X"76",  -- 118
        50708 => X"69",  -- 105
        50709 => X"76",  -- 118
        50710 => X"75",  -- 117
        50711 => X"75",  -- 117
        50712 => X"73",  -- 115
        50713 => X"67",  -- 103
        50714 => X"83",  -- 131
        50715 => X"A1",  -- 161
        50716 => X"9D",  -- 157
        50717 => X"86",  -- 134
        50718 => X"87",  -- 135
        50719 => X"7A",  -- 122
        50720 => X"90",  -- 144
        50721 => X"A6",  -- 166
        50722 => X"AA",  -- 170
        50723 => X"B5",  -- 181
        50724 => X"9A",  -- 154
        50725 => X"A6",  -- 166
        50726 => X"82",  -- 130
        50727 => X"6B",  -- 107
        50728 => X"85",  -- 133
        50729 => X"7E",  -- 126
        50730 => X"2E",  -- 46
        50731 => X"1B",  -- 27
        50732 => X"28",  -- 40
        50733 => X"37",  -- 55
        50734 => X"27",  -- 39
        50735 => X"36",  -- 54
        50736 => X"37",  -- 55
        50737 => X"38",  -- 56
        50738 => X"35",  -- 53
        50739 => X"30",  -- 48
        50740 => X"2F",  -- 47
        50741 => X"32",  -- 50
        50742 => X"31",  -- 49
        50743 => X"2E",  -- 46
        50744 => X"2F",  -- 47
        50745 => X"2C",  -- 44
        50746 => X"2D",  -- 45
        50747 => X"36",  -- 54
        50748 => X"41",  -- 65
        50749 => X"4A",  -- 74
        50750 => X"4A",  -- 74
        50751 => X"46",  -- 70
        50752 => X"43",  -- 67
        50753 => X"43",  -- 67
        50754 => X"40",  -- 64
        50755 => X"3D",  -- 61
        50756 => X"3E",  -- 62
        50757 => X"3F",  -- 63
        50758 => X"3B",  -- 59
        50759 => X"34",  -- 52
        50760 => X"30",  -- 48
        50761 => X"31",  -- 49
        50762 => X"35",  -- 53
        50763 => X"39",  -- 57
        50764 => X"39",  -- 57
        50765 => X"36",  -- 54
        50766 => X"37",  -- 55
        50767 => X"3A",  -- 58
        50768 => X"49",  -- 73
        50769 => X"4A",  -- 74
        50770 => X"49",  -- 73
        50771 => X"44",  -- 68
        50772 => X"43",  -- 67
        50773 => X"47",  -- 71
        50774 => X"4B",  -- 75
        50775 => X"4C",  -- 76
        50776 => X"45",  -- 69
        50777 => X"46",  -- 70
        50778 => X"4A",  -- 74
        50779 => X"48",  -- 72
        50780 => X"49",  -- 73
        50781 => X"61",  -- 97
        50782 => X"82",  -- 130
        50783 => X"94",  -- 148
        50784 => X"85",  -- 133
        50785 => X"78",  -- 120
        50786 => X"7A",  -- 122
        50787 => X"89",  -- 137
        50788 => X"8F",  -- 143
        50789 => X"92",  -- 146
        50790 => X"9D",  -- 157
        50791 => X"A7",  -- 167
        50792 => X"AA",  -- 170
        50793 => X"9A",  -- 154
        50794 => X"92",  -- 146
        50795 => X"9B",  -- 155
        50796 => X"A0",  -- 160
        50797 => X"9F",  -- 159
        50798 => X"9D",  -- 157
        50799 => X"A3",  -- 163
        50800 => X"A9",  -- 169
        50801 => X"A2",  -- 162
        50802 => X"BA",  -- 186
        50803 => X"B9",  -- 185
        50804 => X"B1",  -- 177
        50805 => X"A7",  -- 167
        50806 => X"B4",  -- 180
        50807 => X"A8",  -- 168
        50808 => X"A1",  -- 161
        50809 => X"A7",  -- 167
        50810 => X"A1",  -- 161
        50811 => X"A3",  -- 163
        50812 => X"A2",  -- 162
        50813 => X"A3",  -- 163
        50814 => X"AC",  -- 172
        50815 => X"A7",  -- 167
        50816 => X"A2",  -- 162
        50817 => X"A6",  -- 166
        50818 => X"A8",  -- 168
        50819 => X"A6",  -- 166
        50820 => X"AD",  -- 173
        50821 => X"B7",  -- 183
        50822 => X"BA",  -- 186
        50823 => X"B6",  -- 182
        50824 => X"B9",  -- 185
        50825 => X"B2",  -- 178
        50826 => X"B1",  -- 177
        50827 => X"B8",  -- 184
        50828 => X"BB",  -- 187
        50829 => X"B5",  -- 181
        50830 => X"B2",  -- 178
        50831 => X"B6",  -- 182
        50832 => X"BB",  -- 187
        50833 => X"B7",  -- 183
        50834 => X"B4",  -- 180
        50835 => X"B4",  -- 180
        50836 => X"B6",  -- 182
        50837 => X"B8",  -- 184
        50838 => X"B7",  -- 183
        50839 => X"B6",  -- 182
        50840 => X"B3",  -- 179
        50841 => X"B8",  -- 184
        50842 => X"BB",  -- 187
        50843 => X"BC",  -- 188
        50844 => X"BE",  -- 190
        50845 => X"C3",  -- 195
        50846 => X"C5",  -- 197
        50847 => X"C4",  -- 196
        50848 => X"C7",  -- 199
        50849 => X"C2",  -- 194
        50850 => X"BF",  -- 191
        50851 => X"C0",  -- 192
        50852 => X"C0",  -- 192
        50853 => X"BB",  -- 187
        50854 => X"B7",  -- 183
        50855 => X"B6",  -- 182
        50856 => X"B1",  -- 177
        50857 => X"AE",  -- 174
        50858 => X"A3",  -- 163
        50859 => X"8B",  -- 139
        50860 => X"77",  -- 119
        50861 => X"77",  -- 119
        50862 => X"79",  -- 121
        50863 => X"6D",  -- 109
        50864 => X"56",  -- 86
        50865 => X"46",  -- 70
        50866 => X"39",  -- 57
        50867 => X"31",  -- 49
        50868 => X"2D",  -- 45
        50869 => X"36",  -- 54
        50870 => X"45",  -- 69
        50871 => X"4D",  -- 77
        50872 => X"61",  -- 97
        50873 => X"5D",  -- 93
        50874 => X"65",  -- 101
        50875 => X"77",  -- 119
        50876 => X"8D",  -- 141
        50877 => X"9B",  -- 155
        50878 => X"A5",  -- 165
        50879 => X"AD",  -- 173
        50880 => X"44",  -- 68
        50881 => X"43",  -- 67
        50882 => X"43",  -- 67
        50883 => X"46",  -- 70
        50884 => X"4B",  -- 75
        50885 => X"4D",  -- 77
        50886 => X"4D",  -- 77
        50887 => X"4B",  -- 75
        50888 => X"4E",  -- 78
        50889 => X"46",  -- 70
        50890 => X"40",  -- 64
        50891 => X"41",  -- 65
        50892 => X"49",  -- 73
        50893 => X"51",  -- 81
        50894 => X"51",  -- 81
        50895 => X"50",  -- 80
        50896 => X"47",  -- 71
        50897 => X"45",  -- 69
        50898 => X"44",  -- 68
        50899 => X"43",  -- 67
        50900 => X"43",  -- 67
        50901 => X"42",  -- 66
        50902 => X"40",  -- 64
        50903 => X"3F",  -- 63
        50904 => X"3F",  -- 63
        50905 => X"3D",  -- 61
        50906 => X"3A",  -- 58
        50907 => X"3A",  -- 58
        50908 => X"3C",  -- 60
        50909 => X"3B",  -- 59
        50910 => X"39",  -- 57
        50911 => X"36",  -- 54
        50912 => X"2D",  -- 45
        50913 => X"31",  -- 49
        50914 => X"29",  -- 41
        50915 => X"29",  -- 41
        50916 => X"32",  -- 50
        50917 => X"2E",  -- 46
        50918 => X"2D",  -- 45
        50919 => X"3F",  -- 63
        50920 => X"48",  -- 72
        50921 => X"3F",  -- 63
        50922 => X"39",  -- 57
        50923 => X"34",  -- 52
        50924 => X"51",  -- 81
        50925 => X"5E",  -- 94
        50926 => X"41",  -- 65
        50927 => X"3E",  -- 62
        50928 => X"50",  -- 80
        50929 => X"54",  -- 84
        50930 => X"62",  -- 98
        50931 => X"4F",  -- 79
        50932 => X"4F",  -- 79
        50933 => X"40",  -- 64
        50934 => X"38",  -- 56
        50935 => X"3E",  -- 62
        50936 => X"3A",  -- 58
        50937 => X"30",  -- 48
        50938 => X"38",  -- 56
        50939 => X"66",  -- 102
        50940 => X"6D",  -- 109
        50941 => X"70",  -- 112
        50942 => X"59",  -- 89
        50943 => X"4E",  -- 78
        50944 => X"4C",  -- 76
        50945 => X"42",  -- 66
        50946 => X"4B",  -- 75
        50947 => X"4A",  -- 74
        50948 => X"4A",  -- 74
        50949 => X"52",  -- 82
        50950 => X"49",  -- 73
        50951 => X"43",  -- 67
        50952 => X"32",  -- 50
        50953 => X"3F",  -- 63
        50954 => X"3B",  -- 59
        50955 => X"3D",  -- 61
        50956 => X"4D",  -- 77
        50957 => X"46",  -- 70
        50958 => X"43",  -- 67
        50959 => X"59",  -- 89
        50960 => X"5F",  -- 95
        50961 => X"5A",  -- 90
        50962 => X"5C",  -- 92
        50963 => X"69",  -- 105
        50964 => X"6C",  -- 108
        50965 => X"82",  -- 130
        50966 => X"7F",  -- 127
        50967 => X"8F",  -- 143
        50968 => X"77",  -- 119
        50969 => X"7F",  -- 127
        50970 => X"7D",  -- 125
        50971 => X"7B",  -- 123
        50972 => X"84",  -- 132
        50973 => X"85",  -- 133
        50974 => X"7C",  -- 124
        50975 => X"76",  -- 118
        50976 => X"7D",  -- 125
        50977 => X"5E",  -- 94
        50978 => X"6E",  -- 110
        50979 => X"8F",  -- 143
        50980 => X"85",  -- 133
        50981 => X"82",  -- 130
        50982 => X"86",  -- 134
        50983 => X"7C",  -- 124
        50984 => X"84",  -- 132
        50985 => X"71",  -- 113
        50986 => X"86",  -- 134
        50987 => X"81",  -- 129
        50988 => X"6D",  -- 109
        50989 => X"69",  -- 105
        50990 => X"47",  -- 71
        50991 => X"27",  -- 39
        50992 => X"47",  -- 71
        50993 => X"5D",  -- 93
        50994 => X"75",  -- 117
        50995 => X"7D",  -- 125
        50996 => X"79",  -- 121
        50997 => X"7B",  -- 123
        50998 => X"84",  -- 132
        50999 => X"8A",  -- 138
        51000 => X"8A",  -- 138
        51001 => X"82",  -- 130
        51002 => X"8F",  -- 143
        51003 => X"99",  -- 153
        51004 => X"9A",  -- 154
        51005 => X"B0",  -- 176
        51006 => X"C2",  -- 194
        51007 => X"B7",  -- 183
        51008 => X"C4",  -- 196
        51009 => X"D8",  -- 216
        51010 => X"BD",  -- 189
        51011 => X"BB",  -- 187
        51012 => X"80",  -- 128
        51013 => X"40",  -- 64
        51014 => X"35",  -- 53
        51015 => X"5B",  -- 91
        51016 => X"27",  -- 39
        51017 => X"30",  -- 48
        51018 => X"26",  -- 38
        51019 => X"32",  -- 50
        51020 => X"36",  -- 54
        51021 => X"35",  -- 53
        51022 => X"45",  -- 69
        51023 => X"3C",  -- 60
        51024 => X"42",  -- 66
        51025 => X"63",  -- 99
        51026 => X"62",  -- 98
        51027 => X"87",  -- 135
        51028 => X"74",  -- 116
        51029 => X"7A",  -- 122
        51030 => X"74",  -- 116
        51031 => X"71",  -- 113
        51032 => X"77",  -- 119
        51033 => X"65",  -- 101
        51034 => X"83",  -- 131
        51035 => X"A2",  -- 162
        51036 => X"AA",  -- 170
        51037 => X"86",  -- 134
        51038 => X"8A",  -- 138
        51039 => X"7F",  -- 127
        51040 => X"87",  -- 135
        51041 => X"A0",  -- 160
        51042 => X"AC",  -- 172
        51043 => X"BC",  -- 188
        51044 => X"9D",  -- 157
        51045 => X"A4",  -- 164
        51046 => X"72",  -- 114
        51047 => X"51",  -- 81
        51048 => X"74",  -- 116
        51049 => X"78",  -- 120
        51050 => X"23",  -- 35
        51051 => X"12",  -- 18
        51052 => X"21",  -- 33
        51053 => X"45",  -- 69
        51054 => X"30",  -- 48
        51055 => X"37",  -- 55
        51056 => X"37",  -- 55
        51057 => X"38",  -- 56
        51058 => X"35",  -- 53
        51059 => X"32",  -- 50
        51060 => X"32",  -- 50
        51061 => X"34",  -- 52
        51062 => X"32",  -- 50
        51063 => X"2F",  -- 47
        51064 => X"30",  -- 48
        51065 => X"2D",  -- 45
        51066 => X"2D",  -- 45
        51067 => X"34",  -- 52
        51068 => X"41",  -- 65
        51069 => X"4A",  -- 74
        51070 => X"4B",  -- 75
        51071 => X"46",  -- 70
        51072 => X"43",  -- 67
        51073 => X"43",  -- 67
        51074 => X"41",  -- 65
        51075 => X"3E",  -- 62
        51076 => X"3F",  -- 63
        51077 => X"41",  -- 65
        51078 => X"3C",  -- 60
        51079 => X"34",  -- 52
        51080 => X"2E",  -- 46
        51081 => X"32",  -- 50
        51082 => X"38",  -- 56
        51083 => X"3C",  -- 60
        51084 => X"3A",  -- 58
        51085 => X"37",  -- 55
        51086 => X"38",  -- 56
        51087 => X"3B",  -- 59
        51088 => X"4E",  -- 78
        51089 => X"4D",  -- 77
        51090 => X"4B",  -- 75
        51091 => X"4D",  -- 77
        51092 => X"56",  -- 86
        51093 => X"60",  -- 96
        51094 => X"63",  -- 99
        51095 => X"60",  -- 96
        51096 => X"4B",  -- 75
        51097 => X"4C",  -- 76
        51098 => X"4D",  -- 77
        51099 => X"4A",  -- 74
        51100 => X"4C",  -- 76
        51101 => X"63",  -- 99
        51102 => X"7D",  -- 125
        51103 => X"83",  -- 131
        51104 => X"88",  -- 136
        51105 => X"7B",  -- 123
        51106 => X"81",  -- 129
        51107 => X"8A",  -- 138
        51108 => X"81",  -- 129
        51109 => X"86",  -- 134
        51110 => X"97",  -- 151
        51111 => X"9D",  -- 157
        51112 => X"A9",  -- 169
        51113 => X"9A",  -- 154
        51114 => X"94",  -- 148
        51115 => X"9D",  -- 157
        51116 => X"A0",  -- 160
        51117 => X"98",  -- 152
        51118 => X"9C",  -- 156
        51119 => X"A8",  -- 168
        51120 => X"AD",  -- 173
        51121 => X"99",  -- 153
        51122 => X"B1",  -- 177
        51123 => X"BD",  -- 189
        51124 => X"B6",  -- 182
        51125 => X"A6",  -- 166
        51126 => X"B4",  -- 180
        51127 => X"AD",  -- 173
        51128 => X"A7",  -- 167
        51129 => X"AF",  -- 175
        51130 => X"A1",  -- 161
        51131 => X"9C",  -- 156
        51132 => X"9E",  -- 158
        51133 => X"9C",  -- 156
        51134 => X"A1",  -- 161
        51135 => X"9F",  -- 159
        51136 => X"A3",  -- 163
        51137 => X"A8",  -- 168
        51138 => X"A8",  -- 168
        51139 => X"A1",  -- 161
        51140 => X"A6",  -- 166
        51141 => X"B6",  -- 182
        51142 => X"BD",  -- 189
        51143 => X"B8",  -- 184
        51144 => X"B8",  -- 184
        51145 => X"B5",  -- 181
        51146 => X"B7",  -- 183
        51147 => X"BB",  -- 187
        51148 => X"BB",  -- 187
        51149 => X"B7",  -- 183
        51150 => X"BA",  -- 186
        51151 => X"BF",  -- 191
        51152 => X"BA",  -- 186
        51153 => X"BC",  -- 188
        51154 => X"BC",  -- 188
        51155 => X"B9",  -- 185
        51156 => X"B2",  -- 178
        51157 => X"AD",  -- 173
        51158 => X"AF",  -- 175
        51159 => X"B4",  -- 180
        51160 => X"AC",  -- 172
        51161 => X"B5",  -- 181
        51162 => X"BB",  -- 187
        51163 => X"BA",  -- 186
        51164 => X"BC",  -- 188
        51165 => X"C2",  -- 194
        51166 => X"C6",  -- 198
        51167 => X"C6",  -- 198
        51168 => X"C6",  -- 198
        51169 => X"C0",  -- 192
        51170 => X"BE",  -- 190
        51171 => X"BE",  -- 190
        51172 => X"BE",  -- 190
        51173 => X"B9",  -- 185
        51174 => X"B4",  -- 180
        51175 => X"B2",  -- 178
        51176 => X"AC",  -- 172
        51177 => X"A5",  -- 165
        51178 => X"9D",  -- 157
        51179 => X"8E",  -- 142
        51180 => X"7A",  -- 122
        51181 => X"72",  -- 114
        51182 => X"6F",  -- 111
        51183 => X"66",  -- 102
        51184 => X"4D",  -- 77
        51185 => X"3C",  -- 60
        51186 => X"39",  -- 57
        51187 => X"34",  -- 52
        51188 => X"27",  -- 39
        51189 => X"30",  -- 48
        51190 => X"49",  -- 73
        51191 => X"56",  -- 86
        51192 => X"6D",  -- 109
        51193 => X"71",  -- 113
        51194 => X"75",  -- 117
        51195 => X"7D",  -- 125
        51196 => X"8D",  -- 141
        51197 => X"A0",  -- 160
        51198 => X"AA",  -- 170
        51199 => X"AC",  -- 172
        51200 => X"3B",  -- 59
        51201 => X"3E",  -- 62
        51202 => X"41",  -- 65
        51203 => X"44",  -- 68
        51204 => X"46",  -- 70
        51205 => X"48",  -- 72
        51206 => X"4B",  -- 75
        51207 => X"4D",  -- 77
        51208 => X"53",  -- 83
        51209 => X"45",  -- 69
        51210 => X"3C",  -- 60
        51211 => X"3C",  -- 60
        51212 => X"41",  -- 65
        51213 => X"43",  -- 67
        51214 => X"46",  -- 70
        51215 => X"49",  -- 73
        51216 => X"44",  -- 68
        51217 => X"40",  -- 64
        51218 => X"3D",  -- 61
        51219 => X"3C",  -- 60
        51220 => X"3E",  -- 62
        51221 => X"40",  -- 64
        51222 => X"3E",  -- 62
        51223 => X"3B",  -- 59
        51224 => X"39",  -- 57
        51225 => X"35",  -- 53
        51226 => X"35",  -- 53
        51227 => X"38",  -- 56
        51228 => X"3E",  -- 62
        51229 => X"44",  -- 68
        51230 => X"3F",  -- 63
        51231 => X"33",  -- 51
        51232 => X"38",  -- 56
        51233 => X"2C",  -- 44
        51234 => X"26",  -- 38
        51235 => X"2C",  -- 44
        51236 => X"32",  -- 50
        51237 => X"35",  -- 53
        51238 => X"39",  -- 57
        51239 => X"3E",  -- 62
        51240 => X"42",  -- 66
        51241 => X"34",  -- 52
        51242 => X"3B",  -- 59
        51243 => X"48",  -- 72
        51244 => X"56",  -- 86
        51245 => X"56",  -- 86
        51246 => X"44",  -- 68
        51247 => X"41",  -- 65
        51248 => X"45",  -- 69
        51249 => X"59",  -- 89
        51250 => X"58",  -- 88
        51251 => X"55",  -- 85
        51252 => X"5C",  -- 92
        51253 => X"4B",  -- 75
        51254 => X"3B",  -- 59
        51255 => X"46",  -- 70
        51256 => X"46",  -- 70
        51257 => X"43",  -- 67
        51258 => X"3B",  -- 59
        51259 => X"69",  -- 105
        51260 => X"8B",  -- 139
        51261 => X"71",  -- 113
        51262 => X"5B",  -- 91
        51263 => X"51",  -- 81
        51264 => X"4E",  -- 78
        51265 => X"4C",  -- 76
        51266 => X"44",  -- 68
        51267 => X"53",  -- 83
        51268 => X"56",  -- 86
        51269 => X"4C",  -- 76
        51270 => X"4F",  -- 79
        51271 => X"39",  -- 57
        51272 => X"35",  -- 53
        51273 => X"44",  -- 68
        51274 => X"31",  -- 49
        51275 => X"22",  -- 34
        51276 => X"3A",  -- 58
        51277 => X"4A",  -- 74
        51278 => X"43",  -- 67
        51279 => X"41",  -- 65
        51280 => X"4E",  -- 78
        51281 => X"5F",  -- 95
        51282 => X"5E",  -- 94
        51283 => X"6B",  -- 107
        51284 => X"6F",  -- 111
        51285 => X"6A",  -- 106
        51286 => X"7E",  -- 126
        51287 => X"80",  -- 128
        51288 => X"91",  -- 145
        51289 => X"7D",  -- 125
        51290 => X"73",  -- 115
        51291 => X"7B",  -- 123
        51292 => X"83",  -- 131
        51293 => X"7B",  -- 123
        51294 => X"74",  -- 116
        51295 => X"71",  -- 113
        51296 => X"76",  -- 118
        51297 => X"75",  -- 117
        51298 => X"76",  -- 118
        51299 => X"76",  -- 118
        51300 => X"85",  -- 133
        51301 => X"84",  -- 132
        51302 => X"72",  -- 114
        51303 => X"7E",  -- 126
        51304 => X"8B",  -- 139
        51305 => X"86",  -- 134
        51306 => X"63",  -- 99
        51307 => X"63",  -- 99
        51308 => X"65",  -- 101
        51309 => X"7F",  -- 127
        51310 => X"60",  -- 96
        51311 => X"2A",  -- 42
        51312 => X"4F",  -- 79
        51313 => X"63",  -- 99
        51314 => X"74",  -- 116
        51315 => X"79",  -- 121
        51316 => X"7A",  -- 122
        51317 => X"81",  -- 129
        51318 => X"8D",  -- 141
        51319 => X"95",  -- 149
        51320 => X"93",  -- 147
        51321 => X"8A",  -- 138
        51322 => X"93",  -- 147
        51323 => X"92",  -- 146
        51324 => X"A2",  -- 162
        51325 => X"AD",  -- 173
        51326 => X"C8",  -- 200
        51327 => X"D0",  -- 208
        51328 => X"DF",  -- 223
        51329 => X"DC",  -- 220
        51330 => X"DD",  -- 221
        51331 => X"C3",  -- 195
        51332 => X"8E",  -- 142
        51333 => X"56",  -- 86
        51334 => X"5B",  -- 91
        51335 => X"3F",  -- 63
        51336 => X"48",  -- 72
        51337 => X"3A",  -- 58
        51338 => X"40",  -- 64
        51339 => X"4A",  -- 74
        51340 => X"40",  -- 64
        51341 => X"40",  -- 64
        51342 => X"4C",  -- 76
        51343 => X"4D",  -- 77
        51344 => X"51",  -- 81
        51345 => X"66",  -- 102
        51346 => X"6F",  -- 111
        51347 => X"87",  -- 135
        51348 => X"7B",  -- 123
        51349 => X"7F",  -- 127
        51350 => X"77",  -- 119
        51351 => X"65",  -- 101
        51352 => X"81",  -- 129
        51353 => X"54",  -- 84
        51354 => X"7E",  -- 126
        51355 => X"82",  -- 130
        51356 => X"8C",  -- 140
        51357 => X"A5",  -- 165
        51358 => X"77",  -- 119
        51359 => X"79",  -- 121
        51360 => X"8E",  -- 142
        51361 => X"93",  -- 147
        51362 => X"A9",  -- 169
        51363 => X"BB",  -- 187
        51364 => X"A3",  -- 163
        51365 => X"99",  -- 153
        51366 => X"66",  -- 102
        51367 => X"43",  -- 67
        51368 => X"59",  -- 89
        51369 => X"68",  -- 104
        51370 => X"36",  -- 54
        51371 => X"1A",  -- 26
        51372 => X"2E",  -- 46
        51373 => X"37",  -- 55
        51374 => X"3E",  -- 62
        51375 => X"3D",  -- 61
        51376 => X"3F",  -- 63
        51377 => X"38",  -- 56
        51378 => X"33",  -- 51
        51379 => X"36",  -- 54
        51380 => X"39",  -- 57
        51381 => X"36",  -- 54
        51382 => X"31",  -- 49
        51383 => X"2F",  -- 47
        51384 => X"2C",  -- 44
        51385 => X"2C",  -- 44
        51386 => X"2E",  -- 46
        51387 => X"36",  -- 54
        51388 => X"40",  -- 64
        51389 => X"47",  -- 71
        51390 => X"48",  -- 72
        51391 => X"45",  -- 69
        51392 => X"49",  -- 73
        51393 => X"44",  -- 68
        51394 => X"40",  -- 64
        51395 => X"3F",  -- 63
        51396 => X"40",  -- 64
        51397 => X"3F",  -- 63
        51398 => X"39",  -- 57
        51399 => X"33",  -- 51
        51400 => X"37",  -- 55
        51401 => X"36",  -- 54
        51402 => X"35",  -- 53
        51403 => X"39",  -- 57
        51404 => X"38",  -- 56
        51405 => X"3A",  -- 58
        51406 => X"44",  -- 68
        51407 => X"4F",  -- 79
        51408 => X"57",  -- 87
        51409 => X"5A",  -- 90
        51410 => X"61",  -- 97
        51411 => X"6E",  -- 110
        51412 => X"7E",  -- 126
        51413 => X"84",  -- 132
        51414 => X"7A",  -- 122
        51415 => X"69",  -- 105
        51416 => X"4E",  -- 78
        51417 => X"46",  -- 70
        51418 => X"51",  -- 81
        51419 => X"4D",  -- 77
        51420 => X"4C",  -- 76
        51421 => X"5D",  -- 93
        51422 => X"6F",  -- 111
        51423 => X"83",  -- 131
        51424 => X"83",  -- 131
        51425 => X"7E",  -- 126
        51426 => X"88",  -- 136
        51427 => X"80",  -- 128
        51428 => X"84",  -- 132
        51429 => X"86",  -- 134
        51430 => X"9B",  -- 155
        51431 => X"9B",  -- 155
        51432 => X"A8",  -- 168
        51433 => X"A2",  -- 162
        51434 => X"97",  -- 151
        51435 => X"8D",  -- 141
        51436 => X"92",  -- 146
        51437 => X"A7",  -- 167
        51438 => X"AB",  -- 171
        51439 => X"96",  -- 150
        51440 => X"B2",  -- 178
        51441 => X"97",  -- 151
        51442 => X"9E",  -- 158
        51443 => X"A2",  -- 162
        51444 => X"B3",  -- 179
        51445 => X"B5",  -- 181
        51446 => X"BE",  -- 190
        51447 => X"AE",  -- 174
        51448 => X"B7",  -- 183
        51449 => X"B6",  -- 182
        51450 => X"A0",  -- 160
        51451 => X"AE",  -- 174
        51452 => X"A7",  -- 167
        51453 => X"AA",  -- 170
        51454 => X"A2",  -- 162
        51455 => X"9B",  -- 155
        51456 => X"A0",  -- 160
        51457 => X"A3",  -- 163
        51458 => X"9B",  -- 155
        51459 => X"A5",  -- 165
        51460 => X"AD",  -- 173
        51461 => X"A6",  -- 166
        51462 => X"AF",  -- 175
        51463 => X"BA",  -- 186
        51464 => X"BE",  -- 190
        51465 => X"B2",  -- 178
        51466 => X"B3",  -- 179
        51467 => X"BA",  -- 186
        51468 => X"BB",  -- 187
        51469 => X"BC",  -- 188
        51470 => X"BE",  -- 190
        51471 => X"BB",  -- 187
        51472 => X"BE",  -- 190
        51473 => X"BD",  -- 189
        51474 => X"C1",  -- 193
        51475 => X"C4",  -- 196
        51476 => X"BA",  -- 186
        51477 => X"AC",  -- 172
        51478 => X"AD",  -- 173
        51479 => X"B7",  -- 183
        51480 => X"AD",  -- 173
        51481 => X"AF",  -- 175
        51482 => X"B3",  -- 179
        51483 => X"BC",  -- 188
        51484 => X"C0",  -- 192
        51485 => X"C1",  -- 193
        51486 => X"C1",  -- 193
        51487 => X"C3",  -- 195
        51488 => X"BE",  -- 190
        51489 => X"C1",  -- 193
        51490 => X"BF",  -- 191
        51491 => X"BD",  -- 189
        51492 => X"BC",  -- 188
        51493 => X"B8",  -- 184
        51494 => X"AB",  -- 171
        51495 => X"9E",  -- 158
        51496 => X"A1",  -- 161
        51497 => X"9E",  -- 158
        51498 => X"A4",  -- 164
        51499 => X"91",  -- 145
        51500 => X"6D",  -- 109
        51501 => X"6C",  -- 108
        51502 => X"75",  -- 117
        51503 => X"65",  -- 101
        51504 => X"48",  -- 72
        51505 => X"39",  -- 57
        51506 => X"31",  -- 49
        51507 => X"33",  -- 51
        51508 => X"2F",  -- 47
        51509 => X"2A",  -- 42
        51510 => X"36",  -- 54
        51511 => X"4B",  -- 75
        51512 => X"69",  -- 105
        51513 => X"7D",  -- 125
        51514 => X"8C",  -- 140
        51515 => X"8E",  -- 142
        51516 => X"8A",  -- 138
        51517 => X"92",  -- 146
        51518 => X"A4",  -- 164
        51519 => X"B2",  -- 178
        51520 => X"34",  -- 52
        51521 => X"35",  -- 53
        51522 => X"37",  -- 55
        51523 => X"39",  -- 57
        51524 => X"3B",  -- 59
        51525 => X"3F",  -- 63
        51526 => X"44",  -- 68
        51527 => X"48",  -- 72
        51528 => X"49",  -- 73
        51529 => X"3F",  -- 63
        51530 => X"37",  -- 55
        51531 => X"36",  -- 54
        51532 => X"39",  -- 57
        51533 => X"39",  -- 57
        51534 => X"3A",  -- 58
        51535 => X"3C",  -- 60
        51536 => X"39",  -- 57
        51537 => X"3A",  -- 58
        51538 => X"39",  -- 57
        51539 => X"3A",  -- 58
        51540 => X"3B",  -- 59
        51541 => X"3B",  -- 59
        51542 => X"38",  -- 56
        51543 => X"38",  -- 56
        51544 => X"31",  -- 49
        51545 => X"45",  -- 69
        51546 => X"45",  -- 69
        51547 => X"3A",  -- 58
        51548 => X"40",  -- 64
        51549 => X"43",  -- 67
        51550 => X"41",  -- 65
        51551 => X"47",  -- 71
        51552 => X"36",  -- 54
        51553 => X"38",  -- 56
        51554 => X"3C",  -- 60
        51555 => X"3E",  -- 62
        51556 => X"39",  -- 57
        51557 => X"33",  -- 51
        51558 => X"32",  -- 50
        51559 => X"37",  -- 55
        51560 => X"3C",  -- 60
        51561 => X"2D",  -- 45
        51562 => X"37",  -- 55
        51563 => X"45",  -- 69
        51564 => X"54",  -- 84
        51565 => X"55",  -- 85
        51566 => X"40",  -- 64
        51567 => X"3C",  -- 60
        51568 => X"4C",  -- 76
        51569 => X"5F",  -- 95
        51570 => X"54",  -- 84
        51571 => X"44",  -- 68
        51572 => X"4D",  -- 77
        51573 => X"50",  -- 80
        51574 => X"49",  -- 73
        51575 => X"4C",  -- 76
        51576 => X"43",  -- 67
        51577 => X"3F",  -- 63
        51578 => X"43",  -- 67
        51579 => X"80",  -- 128
        51580 => X"A0",  -- 160
        51581 => X"72",  -- 114
        51582 => X"4F",  -- 79
        51583 => X"49",  -- 73
        51584 => X"48",  -- 72
        51585 => X"47",  -- 71
        51586 => X"41",  -- 65
        51587 => X"58",  -- 88
        51588 => X"6C",  -- 108
        51589 => X"69",  -- 105
        51590 => X"62",  -- 98
        51591 => X"49",  -- 73
        51592 => X"31",  -- 49
        51593 => X"44",  -- 68
        51594 => X"43",  -- 67
        51595 => X"3C",  -- 60
        51596 => X"47",  -- 71
        51597 => X"4B",  -- 75
        51598 => X"45",  -- 69
        51599 => X"46",  -- 70
        51600 => X"43",  -- 67
        51601 => X"55",  -- 85
        51602 => X"59",  -- 89
        51603 => X"67",  -- 103
        51604 => X"6B",  -- 107
        51605 => X"6B",  -- 107
        51606 => X"77",  -- 119
        51607 => X"71",  -- 113
        51608 => X"87",  -- 135
        51609 => X"82",  -- 130
        51610 => X"7C",  -- 124
        51611 => X"7E",  -- 126
        51612 => X"86",  -- 134
        51613 => X"89",  -- 137
        51614 => X"7F",  -- 127
        51615 => X"72",  -- 114
        51616 => X"76",  -- 118
        51617 => X"86",  -- 134
        51618 => X"89",  -- 137
        51619 => X"76",  -- 118
        51620 => X"7B",  -- 123
        51621 => X"85",  -- 133
        51622 => X"7A",  -- 122
        51623 => X"7E",  -- 126
        51624 => X"6E",  -- 110
        51625 => X"74",  -- 116
        51626 => X"7A",  -- 122
        51627 => X"6F",  -- 111
        51628 => X"5F",  -- 95
        51629 => X"78",  -- 120
        51630 => X"62",  -- 98
        51631 => X"56",  -- 86
        51632 => X"67",  -- 103
        51633 => X"66",  -- 102
        51634 => X"67",  -- 103
        51635 => X"6C",  -- 108
        51636 => X"7B",  -- 123
        51637 => X"8A",  -- 138
        51638 => X"8E",  -- 142
        51639 => X"8A",  -- 138
        51640 => X"90",  -- 144
        51641 => X"88",  -- 136
        51642 => X"8F",  -- 143
        51643 => X"92",  -- 146
        51644 => X"A3",  -- 163
        51645 => X"A5",  -- 165
        51646 => X"BF",  -- 191
        51647 => X"D5",  -- 213
        51648 => X"E2",  -- 226
        51649 => X"E3",  -- 227
        51650 => X"E1",  -- 225
        51651 => X"D6",  -- 214
        51652 => X"8E",  -- 142
        51653 => X"55",  -- 85
        51654 => X"53",  -- 83
        51655 => X"4B",  -- 75
        51656 => X"4C",  -- 76
        51657 => X"42",  -- 66
        51658 => X"4B",  -- 75
        51659 => X"57",  -- 87
        51660 => X"50",  -- 80
        51661 => X"50",  -- 80
        51662 => X"59",  -- 89
        51663 => X"5A",  -- 90
        51664 => X"52",  -- 82
        51665 => X"65",  -- 101
        51666 => X"72",  -- 114
        51667 => X"83",  -- 131
        51668 => X"76",  -- 118
        51669 => X"73",  -- 115
        51670 => X"77",  -- 119
        51671 => X"6F",  -- 111
        51672 => X"73",  -- 115
        51673 => X"5B",  -- 91
        51674 => X"70",  -- 112
        51675 => X"7D",  -- 125
        51676 => X"92",  -- 146
        51677 => X"99",  -- 153
        51678 => X"80",  -- 128
        51679 => X"6C",  -- 108
        51680 => X"8E",  -- 142
        51681 => X"9E",  -- 158
        51682 => X"A1",  -- 161
        51683 => X"B6",  -- 182
        51684 => X"A9",  -- 169
        51685 => X"88",  -- 136
        51686 => X"64",  -- 100
        51687 => X"39",  -- 57
        51688 => X"54",  -- 84
        51689 => X"53",  -- 83
        51690 => X"27",  -- 39
        51691 => X"1B",  -- 27
        51692 => X"36",  -- 54
        51693 => X"46",  -- 70
        51694 => X"51",  -- 81
        51695 => X"4D",  -- 77
        51696 => X"44",  -- 68
        51697 => X"3E",  -- 62
        51698 => X"3A",  -- 58
        51699 => X"3B",  -- 59
        51700 => X"3C",  -- 60
        51701 => X"37",  -- 55
        51702 => X"33",  -- 51
        51703 => X"30",  -- 48
        51704 => X"2D",  -- 45
        51705 => X"2C",  -- 44
        51706 => X"30",  -- 48
        51707 => X"36",  -- 54
        51708 => X"3E",  -- 62
        51709 => X"43",  -- 67
        51710 => X"46",  -- 70
        51711 => X"45",  -- 69
        51712 => X"40",  -- 64
        51713 => X"42",  -- 66
        51714 => X"43",  -- 67
        51715 => X"44",  -- 68
        51716 => X"42",  -- 66
        51717 => X"3C",  -- 60
        51718 => X"36",  -- 54
        51719 => X"31",  -- 49
        51720 => X"34",  -- 52
        51721 => X"35",  -- 53
        51722 => X"39",  -- 57
        51723 => X"3F",  -- 63
        51724 => X"43",  -- 67
        51725 => X"49",  -- 73
        51726 => X"53",  -- 83
        51727 => X"5F",  -- 95
        51728 => X"71",  -- 113
        51729 => X"77",  -- 119
        51730 => X"80",  -- 128
        51731 => X"8A",  -- 138
        51732 => X"91",  -- 145
        51733 => X"90",  -- 144
        51734 => X"80",  -- 128
        51735 => X"6F",  -- 111
        51736 => X"52",  -- 82
        51737 => X"47",  -- 71
        51738 => X"48",  -- 72
        51739 => X"48",  -- 72
        51740 => X"55",  -- 85
        51741 => X"68",  -- 104
        51742 => X"6C",  -- 108
        51743 => X"7A",  -- 122
        51744 => X"86",  -- 134
        51745 => X"7F",  -- 127
        51746 => X"87",  -- 135
        51747 => X"7E",  -- 126
        51748 => X"84",  -- 132
        51749 => X"87",  -- 135
        51750 => X"95",  -- 149
        51751 => X"8E",  -- 142
        51752 => X"9E",  -- 158
        51753 => X"98",  -- 152
        51754 => X"92",  -- 146
        51755 => X"8C",  -- 140
        51756 => X"92",  -- 146
        51757 => X"A2",  -- 162
        51758 => X"A5",  -- 165
        51759 => X"94",  -- 148
        51760 => X"A6",  -- 166
        51761 => X"9D",  -- 157
        51762 => X"A4",  -- 164
        51763 => X"A6",  -- 166
        51764 => X"AE",  -- 174
        51765 => X"B5",  -- 181
        51766 => X"B9",  -- 185
        51767 => X"A5",  -- 165
        51768 => X"B4",  -- 180
        51769 => X"BC",  -- 188
        51770 => X"B0",  -- 176
        51771 => X"BC",  -- 188
        51772 => X"AD",  -- 173
        51773 => X"AA",  -- 170
        51774 => X"A5",  -- 165
        51775 => X"A4",  -- 164
        51776 => X"A3",  -- 163
        51777 => X"A8",  -- 168
        51778 => X"9E",  -- 158
        51779 => X"A2",  -- 162
        51780 => X"A9",  -- 169
        51781 => X"A8",  -- 168
        51782 => X"B4",  -- 180
        51783 => X"BE",  -- 190
        51784 => X"BD",  -- 189
        51785 => X"B4",  -- 180
        51786 => X"B4",  -- 180
        51787 => X"BA",  -- 186
        51788 => X"BB",  -- 187
        51789 => X"BE",  -- 190
        51790 => X"C0",  -- 192
        51791 => X"BF",  -- 191
        51792 => X"C3",  -- 195
        51793 => X"C4",  -- 196
        51794 => X"C6",  -- 198
        51795 => X"C6",  -- 198
        51796 => X"B8",  -- 184
        51797 => X"A9",  -- 169
        51798 => X"A8",  -- 168
        51799 => X"B2",  -- 178
        51800 => X"AB",  -- 171
        51801 => X"AC",  -- 172
        51802 => X"B0",  -- 176
        51803 => X"B9",  -- 185
        51804 => X"BE",  -- 190
        51805 => X"BD",  -- 189
        51806 => X"BE",  -- 190
        51807 => X"C2",  -- 194
        51808 => X"C3",  -- 195
        51809 => X"C3",  -- 195
        51810 => X"BF",  -- 191
        51811 => X"BA",  -- 186
        51812 => X"B8",  -- 184
        51813 => X"B6",  -- 182
        51814 => X"AE",  -- 174
        51815 => X"A5",  -- 165
        51816 => X"95",  -- 149
        51817 => X"93",  -- 147
        51818 => X"A3",  -- 163
        51819 => X"A0",  -- 160
        51820 => X"81",  -- 129
        51821 => X"71",  -- 113
        51822 => X"69",  -- 105
        51823 => X"53",  -- 83
        51824 => X"58",  -- 88
        51825 => X"43",  -- 67
        51826 => X"30",  -- 48
        51827 => X"2C",  -- 44
        51828 => X"33",  -- 51
        51829 => X"3D",  -- 61
        51830 => X"45",  -- 69
        51831 => X"4C",  -- 76
        51832 => X"63",  -- 99
        51833 => X"76",  -- 118
        51834 => X"89",  -- 137
        51835 => X"8E",  -- 142
        51836 => X"8F",  -- 143
        51837 => X"96",  -- 150
        51838 => X"A5",  -- 165
        51839 => X"AE",  -- 174
        51840 => X"2F",  -- 47
        51841 => X"2F",  -- 47
        51842 => X"30",  -- 48
        51843 => X"30",  -- 48
        51844 => X"32",  -- 50
        51845 => X"37",  -- 55
        51846 => X"3C",  -- 60
        51847 => X"40",  -- 64
        51848 => X"46",  -- 70
        51849 => X"40",  -- 64
        51850 => X"3C",  -- 60
        51851 => X"3B",  -- 59
        51852 => X"3A",  -- 58
        51853 => X"37",  -- 55
        51854 => X"37",  -- 55
        51855 => X"38",  -- 56
        51856 => X"3C",  -- 60
        51857 => X"3E",  -- 62
        51858 => X"42",  -- 66
        51859 => X"43",  -- 67
        51860 => X"43",  -- 67
        51861 => X"40",  -- 64
        51862 => X"3E",  -- 62
        51863 => X"3E",  -- 62
        51864 => X"4F",  -- 79
        51865 => X"34",  -- 52
        51866 => X"3A",  -- 58
        51867 => X"4B",  -- 75
        51868 => X"48",  -- 72
        51869 => X"49",  -- 73
        51870 => X"4B",  -- 75
        51871 => X"3D",  -- 61
        51872 => X"3A",  -- 58
        51873 => X"4C",  -- 76
        51874 => X"5E",  -- 94
        51875 => X"61",  -- 97
        51876 => X"5B",  -- 91
        51877 => X"5A",  -- 90
        51878 => X"5E",  -- 94
        51879 => X"65",  -- 101
        51880 => X"5A",  -- 90
        51881 => X"59",  -- 89
        51882 => X"63",  -- 99
        51883 => X"61",  -- 97
        51884 => X"54",  -- 84
        51885 => X"49",  -- 73
        51886 => X"3B",  -- 59
        51887 => X"43",  -- 67
        51888 => X"55",  -- 85
        51889 => X"55",  -- 85
        51890 => X"4F",  -- 79
        51891 => X"57",  -- 87
        51892 => X"60",  -- 96
        51893 => X"50",  -- 80
        51894 => X"43",  -- 67
        51895 => X"50",  -- 80
        51896 => X"4F",  -- 79
        51897 => X"46",  -- 70
        51898 => X"42",  -- 66
        51899 => X"6F",  -- 111
        51900 => X"8C",  -- 140
        51901 => X"69",  -- 105
        51902 => X"45",  -- 69
        51903 => X"3B",  -- 59
        51904 => X"46",  -- 70
        51905 => X"51",  -- 81
        51906 => X"51",  -- 81
        51907 => X"63",  -- 99
        51908 => X"74",  -- 116
        51909 => X"67",  -- 103
        51910 => X"50",  -- 80
        51911 => X"38",  -- 56
        51912 => X"35",  -- 53
        51913 => X"3A",  -- 58
        51914 => X"40",  -- 64
        51915 => X"45",  -- 69
        51916 => X"48",  -- 72
        51917 => X"45",  -- 69
        51918 => X"43",  -- 67
        51919 => X"44",  -- 68
        51920 => X"46",  -- 70
        51921 => X"5A",  -- 90
        51922 => X"5F",  -- 95
        51923 => X"68",  -- 104
        51924 => X"6F",  -- 111
        51925 => X"76",  -- 118
        51926 => X"7E",  -- 126
        51927 => X"72",  -- 114
        51928 => X"73",  -- 115
        51929 => X"7A",  -- 122
        51930 => X"77",  -- 119
        51931 => X"71",  -- 113
        51932 => X"7B",  -- 123
        51933 => X"8B",  -- 139
        51934 => X"83",  -- 131
        51935 => X"70",  -- 112
        51936 => X"74",  -- 116
        51937 => X"84",  -- 132
        51938 => X"89",  -- 137
        51939 => X"75",  -- 117
        51940 => X"72",  -- 114
        51941 => X"7C",  -- 124
        51942 => X"7B",  -- 123
        51943 => X"84",  -- 132
        51944 => X"6B",  -- 107
        51945 => X"66",  -- 102
        51946 => X"7E",  -- 126
        51947 => X"71",  -- 113
        51948 => X"68",  -- 104
        51949 => X"7D",  -- 125
        51950 => X"5B",  -- 91
        51951 => X"61",  -- 97
        51952 => X"77",  -- 119
        51953 => X"6D",  -- 109
        51954 => X"64",  -- 100
        51955 => X"6B",  -- 107
        51956 => X"81",  -- 129
        51957 => X"95",  -- 149
        51958 => X"9A",  -- 154
        51959 => X"95",  -- 149
        51960 => X"A0",  -- 160
        51961 => X"96",  -- 150
        51962 => X"93",  -- 147
        51963 => X"8C",  -- 140
        51964 => X"90",  -- 144
        51965 => X"7B",  -- 123
        51966 => X"96",  -- 150
        51967 => X"C5",  -- 197
        51968 => X"E0",  -- 224
        51969 => X"E1",  -- 225
        51970 => X"D7",  -- 215
        51971 => X"CF",  -- 207
        51972 => X"7A",  -- 122
        51973 => X"4A",  -- 74
        51974 => X"47",  -- 71
        51975 => X"56",  -- 86
        51976 => X"61",  -- 97
        51977 => X"5A",  -- 90
        51978 => X"62",  -- 98
        51979 => X"6E",  -- 110
        51980 => X"6C",  -- 108
        51981 => X"6B",  -- 107
        51982 => X"70",  -- 112
        51983 => X"6F",  -- 111
        51984 => X"63",  -- 99
        51985 => X"6C",  -- 108
        51986 => X"7D",  -- 125
        51987 => X"8C",  -- 140
        51988 => X"89",  -- 137
        51989 => X"76",  -- 118
        51990 => X"78",  -- 120
        51991 => X"69",  -- 105
        51992 => X"87",  -- 135
        51993 => X"73",  -- 115
        51994 => X"5E",  -- 94
        51995 => X"6A",  -- 106
        51996 => X"96",  -- 150
        51997 => X"91",  -- 145
        51998 => X"92",  -- 146
        51999 => X"63",  -- 99
        52000 => X"8C",  -- 140
        52001 => X"A8",  -- 168
        52002 => X"9F",  -- 159
        52003 => X"B3",  -- 179
        52004 => X"B9",  -- 185
        52005 => X"81",  -- 129
        52006 => X"63",  -- 99
        52007 => X"36",  -- 54
        52008 => X"50",  -- 80
        52009 => X"3A",  -- 58
        52010 => X"18",  -- 24
        52011 => X"1E",  -- 30
        52012 => X"39",  -- 57
        52013 => X"4C",  -- 76
        52014 => X"55",  -- 85
        52015 => X"4A",  -- 74
        52016 => X"45",  -- 69
        52017 => X"40",  -- 64
        52018 => X"3C",  -- 60
        52019 => X"3E",  -- 62
        52020 => X"3D",  -- 61
        52021 => X"38",  -- 56
        52022 => X"33",  -- 51
        52023 => X"32",  -- 50
        52024 => X"32",  -- 50
        52025 => X"32",  -- 50
        52026 => X"33",  -- 51
        52027 => X"36",  -- 54
        52028 => X"3B",  -- 59
        52029 => X"3E",  -- 62
        52030 => X"42",  -- 66
        52031 => X"44",  -- 68
        52032 => X"3B",  -- 59
        52033 => X"41",  -- 65
        52034 => X"47",  -- 71
        52035 => X"48",  -- 72
        52036 => X"43",  -- 67
        52037 => X"3C",  -- 60
        52038 => X"38",  -- 56
        52039 => X"37",  -- 55
        52040 => X"35",  -- 53
        52041 => X"38",  -- 56
        52042 => X"3C",  -- 60
        52043 => X"43",  -- 67
        52044 => X"4C",  -- 76
        52045 => X"57",  -- 87
        52046 => X"69",  -- 105
        52047 => X"77",  -- 119
        52048 => X"88",  -- 136
        52049 => X"90",  -- 144
        52050 => X"98",  -- 152
        52051 => X"99",  -- 153
        52052 => X"93",  -- 147
        52053 => X"87",  -- 135
        52054 => X"72",  -- 114
        52055 => X"63",  -- 99
        52056 => X"4D",  -- 77
        52057 => X"48",  -- 72
        52058 => X"45",  -- 69
        52059 => X"48",  -- 72
        52060 => X"62",  -- 98
        52061 => X"70",  -- 112
        52062 => X"6E",  -- 110
        52063 => X"7F",  -- 127
        52064 => X"8E",  -- 142
        52065 => X"86",  -- 134
        52066 => X"89",  -- 137
        52067 => X"7D",  -- 125
        52068 => X"88",  -- 136
        52069 => X"8D",  -- 141
        52070 => X"97",  -- 151
        52071 => X"86",  -- 134
        52072 => X"9D",  -- 157
        52073 => X"93",  -- 147
        52074 => X"91",  -- 145
        52075 => X"94",  -- 148
        52076 => X"97",  -- 151
        52077 => X"A1",  -- 161
        52078 => X"A4",  -- 164
        52079 => X"9B",  -- 155
        52080 => X"A0",  -- 160
        52081 => X"A7",  -- 167
        52082 => X"AA",  -- 170
        52083 => X"AA",  -- 170
        52084 => X"A5",  -- 165
        52085 => X"B6",  -- 182
        52086 => X"B5",  -- 181
        52087 => X"A6",  -- 166
        52088 => X"A7",  -- 167
        52089 => X"B6",  -- 182
        52090 => X"B2",  -- 178
        52091 => X"B7",  -- 183
        52092 => X"A7",  -- 167
        52093 => X"A4",  -- 164
        52094 => X"A8",  -- 168
        52095 => X"A9",  -- 169
        52096 => X"9D",  -- 157
        52097 => X"A9",  -- 169
        52098 => X"A1",  -- 161
        52099 => X"A0",  -- 160
        52100 => X"A4",  -- 164
        52101 => X"A3",  -- 163
        52102 => X"AD",  -- 173
        52103 => X"B2",  -- 178
        52104 => X"B9",  -- 185
        52105 => X"B5",  -- 181
        52106 => X"B4",  -- 180
        52107 => X"B9",  -- 185
        52108 => X"BE",  -- 190
        52109 => X"C2",  -- 194
        52110 => X"C3",  -- 195
        52111 => X"C5",  -- 197
        52112 => X"C8",  -- 200
        52113 => X"CA",  -- 202
        52114 => X"CD",  -- 205
        52115 => X"C7",  -- 199
        52116 => X"B5",  -- 181
        52117 => X"A5",  -- 165
        52118 => X"A4",  -- 164
        52119 => X"AC",  -- 172
        52120 => X"AA",  -- 170
        52121 => X"A9",  -- 169
        52122 => X"AC",  -- 172
        52123 => X"B4",  -- 180
        52124 => X"BA",  -- 186
        52125 => X"BA",  -- 186
        52126 => X"BC",  -- 188
        52127 => X"BF",  -- 191
        52128 => X"BE",  -- 190
        52129 => X"BF",  -- 191
        52130 => X"BC",  -- 188
        52131 => X"B8",  -- 184
        52132 => X"B5",  -- 181
        52133 => X"B1",  -- 177
        52134 => X"AB",  -- 171
        52135 => X"A4",  -- 164
        52136 => X"86",  -- 134
        52137 => X"80",  -- 128
        52138 => X"93",  -- 147
        52139 => X"A3",  -- 163
        52140 => X"91",  -- 145
        52141 => X"7C",  -- 124
        52142 => X"6D",  -- 109
        52143 => X"5D",  -- 93
        52144 => X"44",  -- 68
        52145 => X"42",  -- 66
        52146 => X"3D",  -- 61
        52147 => X"37",  -- 55
        52148 => X"39",  -- 57
        52149 => X"42",  -- 66
        52150 => X"4B",  -- 75
        52151 => X"4F",  -- 79
        52152 => X"55",  -- 85
        52153 => X"6C",  -- 108
        52154 => X"88",  -- 136
        52155 => X"99",  -- 153
        52156 => X"A2",  -- 162
        52157 => X"A5",  -- 165
        52158 => X"A8",  -- 168
        52159 => X"A8",  -- 168
        52160 => X"35",  -- 53
        52161 => X"35",  -- 53
        52162 => X"35",  -- 53
        52163 => X"35",  -- 53
        52164 => X"35",  -- 53
        52165 => X"38",  -- 56
        52166 => X"3B",  -- 59
        52167 => X"3E",  -- 62
        52168 => X"48",  -- 72
        52169 => X"47",  -- 71
        52170 => X"46",  -- 70
        52171 => X"45",  -- 69
        52172 => X"44",  -- 68
        52173 => X"42",  -- 66
        52174 => X"41",  -- 65
        52175 => X"41",  -- 65
        52176 => X"49",  -- 73
        52177 => X"4D",  -- 77
        52178 => X"50",  -- 80
        52179 => X"51",  -- 81
        52180 => X"4D",  -- 77
        52181 => X"4A",  -- 74
        52182 => X"48",  -- 72
        52183 => X"49",  -- 73
        52184 => X"3D",  -- 61
        52185 => X"4E",  -- 78
        52186 => X"42",  -- 66
        52187 => X"39",  -- 57
        52188 => X"47",  -- 71
        52189 => X"46",  -- 70
        52190 => X"48",  -- 72
        52191 => X"63",  -- 99
        52192 => X"6E",  -- 110
        52193 => X"7B",  -- 123
        52194 => X"7E",  -- 126
        52195 => X"6F",  -- 111
        52196 => X"5C",  -- 92
        52197 => X"54",  -- 84
        52198 => X"52",  -- 82
        52199 => X"4F",  -- 79
        52200 => X"58",  -- 88
        52201 => X"51",  -- 81
        52202 => X"64",  -- 100
        52203 => X"7D",  -- 125
        52204 => X"94",  -- 148
        52205 => X"93",  -- 147
        52206 => X"6F",  -- 111
        52207 => X"5A",  -- 90
        52208 => X"6C",  -- 108
        52209 => X"5C",  -- 92
        52210 => X"47",  -- 71
        52211 => X"43",  -- 67
        52212 => X"45",  -- 69
        52213 => X"3B",  -- 59
        52214 => X"3E",  -- 62
        52215 => X"54",  -- 84
        52216 => X"44",  -- 68
        52217 => X"35",  -- 53
        52218 => X"3A",  -- 58
        52219 => X"70",  -- 112
        52220 => X"89",  -- 137
        52221 => X"56",  -- 86
        52222 => X"22",  -- 34
        52223 => X"1E",  -- 30
        52224 => X"3D",  -- 61
        52225 => X"51",  -- 81
        52226 => X"5B",  -- 91
        52227 => X"63",  -- 99
        52228 => X"69",  -- 105
        52229 => X"5D",  -- 93
        52230 => X"4D",  -- 77
        52231 => X"47",  -- 71
        52232 => X"42",  -- 66
        52233 => X"31",  -- 49
        52234 => X"2E",  -- 46
        52235 => X"39",  -- 57
        52236 => X"40",  -- 64
        52237 => X"43",  -- 67
        52238 => X"44",  -- 68
        52239 => X"42",  -- 66
        52240 => X"4B",  -- 75
        52241 => X"61",  -- 97
        52242 => X"69",  -- 105
        52243 => X"68",  -- 104
        52244 => X"6C",  -- 108
        52245 => X"79",  -- 121
        52246 => X"82",  -- 130
        52247 => X"7D",  -- 125
        52248 => X"6E",  -- 110
        52249 => X"75",  -- 117
        52250 => X"72",  -- 114
        52251 => X"6B",  -- 107
        52252 => X"75",  -- 117
        52253 => X"87",  -- 135
        52254 => X"84",  -- 132
        52255 => X"74",  -- 116
        52256 => X"7B",  -- 123
        52257 => X"75",  -- 117
        52258 => X"7B",  -- 123
        52259 => X"78",  -- 120
        52260 => X"75",  -- 117
        52261 => X"72",  -- 114
        52262 => X"6F",  -- 111
        52263 => X"82",  -- 130
        52264 => X"79",  -- 121
        52265 => X"6B",  -- 107
        52266 => X"75",  -- 117
        52267 => X"72",  -- 114
        52268 => X"75",  -- 117
        52269 => X"76",  -- 118
        52270 => X"4F",  -- 79
        52271 => X"4D",  -- 77
        52272 => X"6A",  -- 106
        52273 => X"69",  -- 105
        52274 => X"69",  -- 105
        52275 => X"6F",  -- 111
        52276 => X"7A",  -- 122
        52277 => X"88",  -- 136
        52278 => X"95",  -- 149
        52279 => X"9B",  -- 155
        52280 => X"A4",  -- 164
        52281 => X"A1",  -- 161
        52282 => X"98",  -- 152
        52283 => X"84",  -- 132
        52284 => X"74",  -- 116
        52285 => X"4C",  -- 76
        52286 => X"6F",  -- 111
        52287 => X"B9",  -- 185
        52288 => X"EE",  -- 238
        52289 => X"E8",  -- 232
        52290 => X"D8",  -- 216
        52291 => X"BE",  -- 190
        52292 => X"7F",  -- 127
        52293 => X"6A",  -- 106
        52294 => X"80",  -- 128
        52295 => X"9E",  -- 158
        52296 => X"9E",  -- 158
        52297 => X"9A",  -- 154
        52298 => X"9C",  -- 156
        52299 => X"A1",  -- 161
        52300 => X"A0",  -- 160
        52301 => X"9E",  -- 158
        52302 => X"A2",  -- 162
        52303 => X"A3",  -- 163
        52304 => X"9F",  -- 159
        52305 => X"8C",  -- 140
        52306 => X"85",  -- 133
        52307 => X"85",  -- 133
        52308 => X"8C",  -- 140
        52309 => X"77",  -- 119
        52310 => X"7B",  -- 123
        52311 => X"68",  -- 104
        52312 => X"7F",  -- 127
        52313 => X"83",  -- 131
        52314 => X"6E",  -- 110
        52315 => X"61",  -- 97
        52316 => X"83",  -- 131
        52317 => X"71",  -- 113
        52318 => X"8A",  -- 138
        52319 => X"6E",  -- 110
        52320 => X"80",  -- 128
        52321 => X"A0",  -- 160
        52322 => X"A1",  -- 161
        52323 => X"AD",  -- 173
        52324 => X"C4",  -- 196
        52325 => X"85",  -- 133
        52326 => X"5B",  -- 91
        52327 => X"36",  -- 54
        52328 => X"47",  -- 71
        52329 => X"27",  -- 39
        52330 => X"17",  -- 23
        52331 => X"2A",  -- 42
        52332 => X"3D",  -- 61
        52333 => X"4A",  -- 74
        52334 => X"4E",  -- 78
        52335 => X"40",  -- 64
        52336 => X"3F",  -- 63
        52337 => X"3B",  -- 59
        52338 => X"3B",  -- 59
        52339 => X"3D",  -- 61
        52340 => X"3B",  -- 59
        52341 => X"37",  -- 55
        52342 => X"34",  -- 52
        52343 => X"35",  -- 53
        52344 => X"3C",  -- 60
        52345 => X"3D",  -- 61
        52346 => X"3B",  -- 59
        52347 => X"3B",  -- 59
        52348 => X"3A",  -- 58
        52349 => X"3B",  -- 59
        52350 => X"3D",  -- 61
        52351 => X"40",  -- 64
        52352 => X"3C",  -- 60
        52353 => X"40",  -- 64
        52354 => X"45",  -- 69
        52355 => X"45",  -- 69
        52356 => X"41",  -- 65
        52357 => X"3D",  -- 61
        52358 => X"3C",  -- 60
        52359 => X"3C",  -- 60
        52360 => X"3B",  -- 59
        52361 => X"3C",  -- 60
        52362 => X"41",  -- 65
        52363 => X"47",  -- 71
        52364 => X"52",  -- 82
        52365 => X"65",  -- 101
        52366 => X"7B",  -- 123
        52367 => X"8B",  -- 139
        52368 => X"95",  -- 149
        52369 => X"97",  -- 151
        52370 => X"97",  -- 151
        52371 => X"8C",  -- 140
        52372 => X"7B",  -- 123
        52373 => X"67",  -- 103
        52374 => X"56",  -- 86
        52375 => X"4C",  -- 76
        52376 => X"44",  -- 68
        52377 => X"4A",  -- 74
        52378 => X"4B",  -- 75
        52379 => X"50",  -- 80
        52380 => X"6B",  -- 107
        52381 => X"76",  -- 118
        52382 => X"73",  -- 115
        52383 => X"92",  -- 146
        52384 => X"90",  -- 144
        52385 => X"87",  -- 135
        52386 => X"88",  -- 136
        52387 => X"79",  -- 121
        52388 => X"82",  -- 130
        52389 => X"8B",  -- 139
        52390 => X"97",  -- 151
        52391 => X"86",  -- 134
        52392 => X"9C",  -- 156
        52393 => X"92",  -- 146
        52394 => X"93",  -- 147
        52395 => X"99",  -- 153
        52396 => X"9A",  -- 154
        52397 => X"9C",  -- 156
        52398 => X"A0",  -- 160
        52399 => X"9E",  -- 158
        52400 => X"9F",  -- 159
        52401 => X"AA",  -- 170
        52402 => X"A6",  -- 166
        52403 => X"A8",  -- 168
        52404 => X"9A",  -- 154
        52405 => X"AE",  -- 174
        52406 => X"AE",  -- 174
        52407 => X"B1",  -- 177
        52408 => X"9D",  -- 157
        52409 => X"AB",  -- 171
        52410 => X"A6",  -- 166
        52411 => X"A5",  -- 165
        52412 => X"9F",  -- 159
        52413 => X"9E",  -- 158
        52414 => X"A9",  -- 169
        52415 => X"A8",  -- 168
        52416 => X"96",  -- 150
        52417 => X"A9",  -- 169
        52418 => X"A6",  -- 166
        52419 => X"A3",  -- 163
        52420 => X"A4",  -- 164
        52421 => X"A0",  -- 160
        52422 => X"A2",  -- 162
        52423 => X"A0",  -- 160
        52424 => X"B1",  -- 177
        52425 => X"B3",  -- 179
        52426 => X"B2",  -- 178
        52427 => X"B6",  -- 182
        52428 => X"BF",  -- 191
        52429 => X"C4",  -- 196
        52430 => X"C5",  -- 197
        52431 => X"C9",  -- 201
        52432 => X"CB",  -- 203
        52433 => X"CF",  -- 207
        52434 => X"D0",  -- 208
        52435 => X"C5",  -- 197
        52436 => X"B1",  -- 177
        52437 => X"A3",  -- 163
        52438 => X"A2",  -- 162
        52439 => X"A8",  -- 168
        52440 => X"AA",  -- 170
        52441 => X"A7",  -- 167
        52442 => X"A9",  -- 169
        52443 => X"AF",  -- 175
        52444 => X"B6",  -- 182
        52445 => X"B7",  -- 183
        52446 => X"B9",  -- 185
        52447 => X"BC",  -- 188
        52448 => X"B3",  -- 179
        52449 => X"B6",  -- 182
        52450 => X"B8",  -- 184
        52451 => X"B8",  -- 184
        52452 => X"B4",  -- 180
        52453 => X"AC",  -- 172
        52454 => X"A2",  -- 162
        52455 => X"9B",  -- 155
        52456 => X"89",  -- 137
        52457 => X"76",  -- 118
        52458 => X"7D",  -- 125
        52459 => X"92",  -- 146
        52460 => X"8F",  -- 143
        52461 => X"7F",  -- 127
        52462 => X"77",  -- 119
        52463 => X"73",  -- 115
        52464 => X"3A",  -- 58
        52465 => X"3C",  -- 60
        52466 => X"3F",  -- 63
        52467 => X"3F",  -- 63
        52468 => X"40",  -- 64
        52469 => X"45",  -- 69
        52470 => X"4F",  -- 79
        52471 => X"59",  -- 89
        52472 => X"55",  -- 85
        52473 => X"64",  -- 100
        52474 => X"7D",  -- 125
        52475 => X"93",  -- 147
        52476 => X"A3",  -- 163
        52477 => X"AB",  -- 171
        52478 => X"AD",  -- 173
        52479 => X"AC",  -- 172
        52480 => X"40",  -- 64
        52481 => X"41",  -- 65
        52482 => X"42",  -- 66
        52483 => X"44",  -- 68
        52484 => X"44",  -- 68
        52485 => X"45",  -- 69
        52486 => X"48",  -- 72
        52487 => X"49",  -- 73
        52488 => X"4F",  -- 79
        52489 => X"4F",  -- 79
        52490 => X"50",  -- 80
        52491 => X"4E",  -- 78
        52492 => X"4D",  -- 77
        52493 => X"4D",  -- 77
        52494 => X"4C",  -- 76
        52495 => X"4B",  -- 75
        52496 => X"4F",  -- 79
        52497 => X"51",  -- 81
        52498 => X"53",  -- 83
        52499 => X"51",  -- 81
        52500 => X"4D",  -- 77
        52501 => X"49",  -- 73
        52502 => X"4A",  -- 74
        52503 => X"4A",  -- 74
        52504 => X"46",  -- 70
        52505 => X"41",  -- 65
        52506 => X"41",  -- 65
        52507 => X"35",  -- 53
        52508 => X"31",  -- 49
        52509 => X"5C",  -- 92
        52510 => X"76",  -- 118
        52511 => X"5C",  -- 92
        52512 => X"31",  -- 49
        52513 => X"39",  -- 57
        52514 => X"3B",  -- 59
        52515 => X"38",  -- 56
        52516 => X"36",  -- 54
        52517 => X"3C",  -- 60
        52518 => X"3E",  -- 62
        52519 => X"3B",  -- 59
        52520 => X"33",  -- 51
        52521 => X"31",  -- 49
        52522 => X"38",  -- 56
        52523 => X"30",  -- 48
        52524 => X"2A",  -- 42
        52525 => X"36",  -- 54
        52526 => X"44",  -- 68
        52527 => X"5C",  -- 92
        52528 => X"87",  -- 135
        52529 => X"98",  -- 152
        52530 => X"8F",  -- 143
        52531 => X"71",  -- 113
        52532 => X"66",  -- 102
        52533 => X"66",  -- 102
        52534 => X"59",  -- 89
        52535 => X"46",  -- 70
        52536 => X"4B",  -- 75
        52537 => X"31",  -- 49
        52538 => X"3E",  -- 62
        52539 => X"74",  -- 116
        52540 => X"78",  -- 120
        52541 => X"32",  -- 50
        52542 => X"09",  -- 9
        52543 => X"25",  -- 37
        52544 => X"46",  -- 70
        52545 => X"54",  -- 84
        52546 => X"60",  -- 96
        52547 => X"5F",  -- 95
        52548 => X"5B",  -- 91
        52549 => X"58",  -- 88
        52550 => X"50",  -- 80
        52551 => X"50",  -- 80
        52552 => X"40",  -- 64
        52553 => X"31",  -- 49
        52554 => X"2F",  -- 47
        52555 => X"39",  -- 57
        52556 => X"3F",  -- 63
        52557 => X"44",  -- 68
        52558 => X"45",  -- 69
        52559 => X"41",  -- 65
        52560 => X"41",  -- 65
        52561 => X"57",  -- 87
        52562 => X"68",  -- 104
        52563 => X"62",  -- 98
        52564 => X"62",  -- 98
        52565 => X"6F",  -- 111
        52566 => X"79",  -- 121
        52567 => X"7B",  -- 123
        52568 => X"7A",  -- 122
        52569 => X"7A",  -- 122
        52570 => X"7B",  -- 123
        52571 => X"7B",  -- 123
        52572 => X"81",  -- 129
        52573 => X"87",  -- 135
        52574 => X"82",  -- 130
        52575 => X"79",  -- 121
        52576 => X"85",  -- 133
        52577 => X"75",  -- 117
        52578 => X"7A",  -- 122
        52579 => X"7D",  -- 125
        52580 => X"7B",  -- 123
        52581 => X"78",  -- 120
        52582 => X"6E",  -- 110
        52583 => X"75",  -- 117
        52584 => X"73",  -- 115
        52585 => X"74",  -- 116
        52586 => X"71",  -- 113
        52587 => X"73",  -- 115
        52588 => X"76",  -- 118
        52589 => X"5D",  -- 93
        52590 => X"50",  -- 80
        52591 => X"55",  -- 85
        52592 => X"65",  -- 101
        52593 => X"6D",  -- 109
        52594 => X"74",  -- 116
        52595 => X"7A",  -- 122
        52596 => X"7E",  -- 126
        52597 => X"86",  -- 134
        52598 => X"91",  -- 145
        52599 => X"9A",  -- 154
        52600 => X"9F",  -- 159
        52601 => X"A8",  -- 168
        52602 => X"A9",  -- 169
        52603 => X"88",  -- 136
        52604 => X"5F",  -- 95
        52605 => X"21",  -- 33
        52606 => X"41",  -- 65
        52607 => X"95",  -- 149
        52608 => X"B7",  -- 183
        52609 => X"D0",  -- 208
        52610 => X"EC",  -- 236
        52611 => X"CF",  -- 207
        52612 => X"A8",  -- 168
        52613 => X"85",  -- 133
        52614 => X"7B",  -- 123
        52615 => X"71",  -- 113
        52616 => X"66",  -- 102
        52617 => X"65",  -- 101
        52618 => X"62",  -- 98
        52619 => X"5F",  -- 95
        52620 => X"5E",  -- 94
        52621 => X"5D",  -- 93
        52622 => X"5E",  -- 94
        52623 => X"66",  -- 102
        52624 => X"77",  -- 119
        52625 => X"73",  -- 115
        52626 => X"84",  -- 132
        52627 => X"9B",  -- 155
        52628 => X"AD",  -- 173
        52629 => X"92",  -- 146
        52630 => X"86",  -- 134
        52631 => X"64",  -- 100
        52632 => X"7F",  -- 127
        52633 => X"7F",  -- 127
        52634 => X"6C",  -- 108
        52635 => X"50",  -- 80
        52636 => X"79",  -- 121
        52637 => X"6C",  -- 108
        52638 => X"6E",  -- 110
        52639 => X"5B",  -- 91
        52640 => X"6F",  -- 111
        52641 => X"8D",  -- 141
        52642 => X"A1",  -- 161
        52643 => X"A3",  -- 163
        52644 => X"BE",  -- 190
        52645 => X"8B",  -- 139
        52646 => X"4A",  -- 74
        52647 => X"2E",  -- 46
        52648 => X"38",  -- 56
        52649 => X"1A",  -- 26
        52650 => X"20",  -- 32
        52651 => X"3A",  -- 58
        52652 => X"43",  -- 67
        52653 => X"46",  -- 70
        52654 => X"44",  -- 68
        52655 => X"3A",  -- 58
        52656 => X"36",  -- 54
        52657 => X"35",  -- 53
        52658 => X"38",  -- 56
        52659 => X"3A",  -- 58
        52660 => X"3B",  -- 59
        52661 => X"38",  -- 56
        52662 => X"39",  -- 57
        52663 => X"3C",  -- 60
        52664 => X"47",  -- 71
        52665 => X"45",  -- 69
        52666 => X"42",  -- 66
        52667 => X"3D",  -- 61
        52668 => X"3A",  -- 58
        52669 => X"38",  -- 56
        52670 => X"3A",  -- 58
        52671 => X"3C",  -- 60
        52672 => X"3E",  -- 62
        52673 => X"41",  -- 65
        52674 => X"45",  -- 69
        52675 => X"46",  -- 70
        52676 => X"43",  -- 67
        52677 => X"3F",  -- 63
        52678 => X"3B",  -- 59
        52679 => X"39",  -- 57
        52680 => X"3C",  -- 60
        52681 => X"44",  -- 68
        52682 => X"4D",  -- 77
        52683 => X"55",  -- 85
        52684 => X"62",  -- 98
        52685 => X"73",  -- 115
        52686 => X"84",  -- 132
        52687 => X"90",  -- 144
        52688 => X"94",  -- 148
        52689 => X"8F",  -- 143
        52690 => X"83",  -- 131
        52691 => X"72",  -- 114
        52692 => X"5E",  -- 94
        52693 => X"4D",  -- 77
        52694 => X"46",  -- 70
        52695 => X"45",  -- 69
        52696 => X"45",  -- 69
        52697 => X"49",  -- 73
        52698 => X"4D",  -- 77
        52699 => X"54",  -- 84
        52700 => X"72",  -- 114
        52701 => X"7C",  -- 124
        52702 => X"79",  -- 121
        52703 => X"98",  -- 152
        52704 => X"8A",  -- 138
        52705 => X"84",  -- 132
        52706 => X"84",  -- 132
        52707 => X"74",  -- 116
        52708 => X"7B",  -- 123
        52709 => X"84",  -- 132
        52710 => X"96",  -- 150
        52711 => X"8C",  -- 140
        52712 => X"93",  -- 147
        52713 => X"88",  -- 136
        52714 => X"8D",  -- 141
        52715 => X"96",  -- 150
        52716 => X"95",  -- 149
        52717 => X"92",  -- 146
        52718 => X"99",  -- 153
        52719 => X"9E",  -- 158
        52720 => X"9C",  -- 156
        52721 => X"A6",  -- 166
        52722 => X"A0",  -- 160
        52723 => X"A7",  -- 167
        52724 => X"9B",  -- 155
        52725 => X"A5",  -- 165
        52726 => X"A6",  -- 166
        52727 => X"B7",  -- 183
        52728 => X"A4",  -- 164
        52729 => X"AC",  -- 172
        52730 => X"A3",  -- 163
        52731 => X"9F",  -- 159
        52732 => X"A2",  -- 162
        52733 => X"A3",  -- 163
        52734 => X"A8",  -- 168
        52735 => X"9A",  -- 154
        52736 => X"97",  -- 151
        52737 => X"AA",  -- 170
        52738 => X"A5",  -- 165
        52739 => X"A3",  -- 163
        52740 => X"A5",  -- 165
        52741 => X"A2",  -- 162
        52742 => X"A4",  -- 164
        52743 => X"A0",  -- 160
        52744 => X"AA",  -- 170
        52745 => X"B3",  -- 179
        52746 => X"B0",  -- 176
        52747 => X"B2",  -- 178
        52748 => X"C0",  -- 192
        52749 => X"C5",  -- 197
        52750 => X"C6",  -- 198
        52751 => X"CE",  -- 206
        52752 => X"CD",  -- 205
        52753 => X"D2",  -- 210
        52754 => X"CF",  -- 207
        52755 => X"BE",  -- 190
        52756 => X"AC",  -- 172
        52757 => X"A1",  -- 161
        52758 => X"A2",  -- 162
        52759 => X"A6",  -- 166
        52760 => X"AC",  -- 172
        52761 => X"A6",  -- 166
        52762 => X"A7",  -- 167
        52763 => X"AC",  -- 172
        52764 => X"B3",  -- 179
        52765 => X"B4",  -- 180
        52766 => X"B6",  -- 182
        52767 => X"B8",  -- 184
        52768 => X"AE",  -- 174
        52769 => X"AF",  -- 175
        52770 => X"B1",  -- 177
        52771 => X"B3",  -- 179
        52772 => X"B1",  -- 177
        52773 => X"A7",  -- 167
        52774 => X"9C",  -- 156
        52775 => X"94",  -- 148
        52776 => X"93",  -- 147
        52777 => X"79",  -- 121
        52778 => X"72",  -- 114
        52779 => X"81",  -- 129
        52780 => X"83",  -- 131
        52781 => X"77",  -- 119
        52782 => X"6F",  -- 111
        52783 => X"6E",  -- 110
        52784 => X"56",  -- 86
        52785 => X"3F",  -- 63
        52786 => X"30",  -- 48
        52787 => X"39",  -- 57
        52788 => X"47",  -- 71
        52789 => X"50",  -- 80
        52790 => X"5B",  -- 91
        52791 => X"67",  -- 103
        52792 => X"65",  -- 101
        52793 => X"68",  -- 104
        52794 => X"70",  -- 112
        52795 => X"7F",  -- 127
        52796 => X"91",  -- 145
        52797 => X"A1",  -- 161
        52798 => X"AC",  -- 172
        52799 => X"B2",  -- 178
        52800 => X"4A",  -- 74
        52801 => X"4C",  -- 76
        52802 => X"4E",  -- 78
        52803 => X"50",  -- 80
        52804 => X"51",  -- 81
        52805 => X"53",  -- 83
        52806 => X"55",  -- 85
        52807 => X"56",  -- 86
        52808 => X"59",  -- 89
        52809 => X"58",  -- 88
        52810 => X"55",  -- 85
        52811 => X"51",  -- 81
        52812 => X"51",  -- 81
        52813 => X"54",  -- 84
        52814 => X"54",  -- 84
        52815 => X"51",  -- 81
        52816 => X"4E",  -- 78
        52817 => X"4F",  -- 79
        52818 => X"4F",  -- 79
        52819 => X"4D",  -- 77
        52820 => X"4A",  -- 74
        52821 => X"46",  -- 70
        52822 => X"46",  -- 70
        52823 => X"44",  -- 68
        52824 => X"48",  -- 72
        52825 => X"3F",  -- 63
        52826 => X"29",  -- 41
        52827 => X"35",  -- 53
        52828 => X"63",  -- 99
        52829 => X"66",  -- 102
        52830 => X"49",  -- 73
        52831 => X"3F",  -- 63
        52832 => X"33",  -- 51
        52833 => X"36",  -- 54
        52834 => X"36",  -- 54
        52835 => X"37",  -- 55
        52836 => X"3A",  -- 58
        52837 => X"3C",  -- 60
        52838 => X"3B",  -- 59
        52839 => X"36",  -- 54
        52840 => X"4D",  -- 77
        52841 => X"45",  -- 69
        52842 => X"45",  -- 69
        52843 => X"3A",  -- 58
        52844 => X"32",  -- 50
        52845 => X"32",  -- 50
        52846 => X"29",  -- 41
        52847 => X"2F",  -- 47
        52848 => X"37",  -- 55
        52849 => X"44",  -- 68
        52850 => X"49",  -- 73
        52851 => X"43",  -- 67
        52852 => X"55",  -- 85
        52853 => X"7B",  -- 123
        52854 => X"94",  -- 148
        52855 => X"98",  -- 152
        52856 => X"59",  -- 89
        52857 => X"5A",  -- 90
        52858 => X"60",  -- 96
        52859 => X"5C",  -- 92
        52860 => X"4C",  -- 76
        52861 => X"26",  -- 38
        52862 => X"11",  -- 17
        52863 => X"2E",  -- 46
        52864 => X"38",  -- 56
        52865 => X"3E",  -- 62
        52866 => X"5A",  -- 90
        52867 => X"5E",  -- 94
        52868 => X"58",  -- 88
        52869 => X"58",  -- 88
        52870 => X"47",  -- 71
        52871 => X"36",  -- 54
        52872 => X"31",  -- 49
        52873 => X"38",  -- 56
        52874 => X"3D",  -- 61
        52875 => X"3E",  -- 62
        52876 => X"40",  -- 64
        52877 => X"40",  -- 64
        52878 => X"3F",  -- 63
        52879 => X"3C",  -- 60
        52880 => X"39",  -- 57
        52881 => X"50",  -- 80
        52882 => X"6C",  -- 108
        52883 => X"66",  -- 102
        52884 => X"61",  -- 97
        52885 => X"6C",  -- 108
        52886 => X"6D",  -- 109
        52887 => X"74",  -- 116
        52888 => X"7B",  -- 123
        52889 => X"7A",  -- 122
        52890 => X"7D",  -- 125
        52891 => X"84",  -- 132
        52892 => X"86",  -- 134
        52893 => X"7F",  -- 127
        52894 => X"74",  -- 116
        52895 => X"6E",  -- 110
        52896 => X"7C",  -- 124
        52897 => X"75",  -- 117
        52898 => X"7F",  -- 127
        52899 => X"7D",  -- 125
        52900 => X"7D",  -- 125
        52901 => X"87",  -- 135
        52902 => X"7E",  -- 126
        52903 => X"71",  -- 113
        52904 => X"69",  -- 105
        52905 => X"6B",  -- 107
        52906 => X"61",  -- 97
        52907 => X"68",  -- 104
        52908 => X"79",  -- 121
        52909 => X"5F",  -- 95
        52910 => X"61",  -- 97
        52911 => X"6B",  -- 107
        52912 => X"65",  -- 101
        52913 => X"69",  -- 105
        52914 => X"70",  -- 112
        52915 => X"7E",  -- 126
        52916 => X"89",  -- 137
        52917 => X"8F",  -- 143
        52918 => X"91",  -- 145
        52919 => X"94",  -- 148
        52920 => X"77",  -- 119
        52921 => X"8F",  -- 143
        52922 => X"A6",  -- 166
        52923 => X"8D",  -- 141
        52924 => X"59",  -- 89
        52925 => X"18",  -- 24
        52926 => X"32",  -- 50
        52927 => X"76",  -- 118
        52928 => X"91",  -- 145
        52929 => X"B3",  -- 179
        52930 => X"D2",  -- 210
        52931 => X"A2",  -- 162
        52932 => X"8E",  -- 142
        52933 => X"86",  -- 134
        52934 => X"8F",  -- 143
        52935 => X"8C",  -- 140
        52936 => X"6D",  -- 109
        52937 => X"73",  -- 115
        52938 => X"70",  -- 112
        52939 => X"69",  -- 105
        52940 => X"68",  -- 104
        52941 => X"64",  -- 100
        52942 => X"65",  -- 101
        52943 => X"71",  -- 113
        52944 => X"6A",  -- 106
        52945 => X"67",  -- 103
        52946 => X"6B",  -- 107
        52947 => X"7A",  -- 122
        52948 => X"86",  -- 134
        52949 => X"85",  -- 133
        52950 => X"94",  -- 148
        52951 => X"8A",  -- 138
        52952 => X"97",  -- 151
        52953 => X"93",  -- 147
        52954 => X"77",  -- 119
        52955 => X"50",  -- 80
        52956 => X"72",  -- 114
        52957 => X"69",  -- 105
        52958 => X"58",  -- 88
        52959 => X"58",  -- 88
        52960 => X"66",  -- 102
        52961 => X"84",  -- 132
        52962 => X"9B",  -- 155
        52963 => X"99",  -- 153
        52964 => X"AE",  -- 174
        52965 => X"8B",  -- 139
        52966 => X"3F",  -- 63
        52967 => X"23",  -- 35
        52968 => X"2B",  -- 43
        52969 => X"16",  -- 22
        52970 => X"29",  -- 41
        52971 => X"3F",  -- 63
        52972 => X"3D",  -- 61
        52973 => X"39",  -- 57
        52974 => X"30",  -- 48
        52975 => X"2F",  -- 47
        52976 => X"33",  -- 51
        52977 => X"33",  -- 51
        52978 => X"37",  -- 55
        52979 => X"3B",  -- 59
        52980 => X"3B",  -- 59
        52981 => X"3A",  -- 58
        52982 => X"3C",  -- 60
        52983 => X"42",  -- 66
        52984 => X"4A",  -- 74
        52985 => X"47",  -- 71
        52986 => X"43",  -- 67
        52987 => X"3D",  -- 61
        52988 => X"3A",  -- 58
        52989 => X"39",  -- 57
        52990 => X"39",  -- 57
        52991 => X"39",  -- 57
        52992 => X"3B",  -- 59
        52993 => X"40",  -- 64
        52994 => X"46",  -- 70
        52995 => X"48",  -- 72
        52996 => X"43",  -- 67
        52997 => X"3D",  -- 61
        52998 => X"37",  -- 55
        52999 => X"34",  -- 52
        53000 => X"41",  -- 65
        53001 => X"4F",  -- 79
        53002 => X"5D",  -- 93
        53003 => X"68",  -- 104
        53004 => X"72",  -- 114
        53005 => X"7B",  -- 123
        53006 => X"83",  -- 131
        53007 => X"86",  -- 134
        53008 => X"82",  -- 130
        53009 => X"77",  -- 119
        53010 => X"67",  -- 103
        53011 => X"58",  -- 88
        53012 => X"4B",  -- 75
        53013 => X"42",  -- 66
        53014 => X"43",  -- 67
        53015 => X"48",  -- 72
        53016 => X"4F",  -- 79
        53017 => X"47",  -- 71
        53018 => X"49",  -- 73
        53019 => X"58",  -- 88
        53020 => X"78",  -- 120
        53021 => X"84",  -- 132
        53022 => X"7D",  -- 125
        53023 => X"8F",  -- 143
        53024 => X"8E",  -- 142
        53025 => X"86",  -- 134
        53026 => X"8A",  -- 138
        53027 => X"7E",  -- 126
        53028 => X"82",  -- 130
        53029 => X"86",  -- 134
        53030 => X"98",  -- 152
        53031 => X"94",  -- 148
        53032 => X"89",  -- 137
        53033 => X"85",  -- 133
        53034 => X"8D",  -- 141
        53035 => X"97",  -- 151
        53036 => X"93",  -- 147
        53037 => X"90",  -- 144
        53038 => X"99",  -- 153
        53039 => X"9E",  -- 158
        53040 => X"98",  -- 152
        53041 => X"A1",  -- 161
        53042 => X"A1",  -- 161
        53043 => X"A9",  -- 169
        53044 => X"A6",  -- 166
        53045 => X"A5",  -- 165
        53046 => X"A3",  -- 163
        53047 => X"B5",  -- 181
        53048 => X"AE",  -- 174
        53049 => X"B2",  -- 178
        53050 => X"AA",  -- 170
        53051 => X"A0",  -- 160
        53052 => X"AA",  -- 170
        53053 => X"A4",  -- 164
        53054 => X"A2",  -- 162
        53055 => X"87",  -- 135
        53056 => X"99",  -- 153
        53057 => X"A5",  -- 165
        53058 => X"9A",  -- 154
        53059 => X"9C",  -- 156
        53060 => X"A3",  -- 163
        53061 => X"A2",  -- 162
        53062 => X"AB",  -- 171
        53063 => X"AC",  -- 172
        53064 => X"A8",  -- 168
        53065 => X"B6",  -- 182
        53066 => X"B1",  -- 177
        53067 => X"B0",  -- 176
        53068 => X"C0",  -- 192
        53069 => X"C5",  -- 197
        53070 => X"C4",  -- 196
        53071 => X"CD",  -- 205
        53072 => X"CF",  -- 207
        53073 => X"D1",  -- 209
        53074 => X"C9",  -- 201
        53075 => X"B6",  -- 182
        53076 => X"A3",  -- 163
        53077 => X"9F",  -- 159
        53078 => X"A3",  -- 163
        53079 => X"A4",  -- 164
        53080 => X"AD",  -- 173
        53081 => X"A6",  -- 166
        53082 => X"A6",  -- 166
        53083 => X"AA",  -- 170
        53084 => X"B0",  -- 176
        53085 => X"B0",  -- 176
        53086 => X"B0",  -- 176
        53087 => X"B1",  -- 177
        53088 => X"B3",  -- 179
        53089 => X"AD",  -- 173
        53090 => X"A9",  -- 169
        53091 => X"AA",  -- 170
        53092 => X"A9",  -- 169
        53093 => X"A1",  -- 161
        53094 => X"97",  -- 151
        53095 => X"91",  -- 145
        53096 => X"8B",  -- 139
        53097 => X"78",  -- 120
        53098 => X"6C",  -- 108
        53099 => X"73",  -- 115
        53100 => X"7A",  -- 122
        53101 => X"70",  -- 112
        53102 => X"63",  -- 99
        53103 => X"5C",  -- 92
        53104 => X"57",  -- 87
        53105 => X"41",  -- 65
        53106 => X"36",  -- 54
        53107 => X"42",  -- 66
        53108 => X"4C",  -- 76
        53109 => X"4F",  -- 79
        53110 => X"5B",  -- 91
        53111 => X"6C",  -- 108
        53112 => X"70",  -- 112
        53113 => X"6E",  -- 110
        53114 => X"73",  -- 115
        53115 => X"80",  -- 128
        53116 => X"90",  -- 144
        53117 => X"9C",  -- 156
        53118 => X"A3",  -- 163
        53119 => X"A8",  -- 168
        53120 => X"4E",  -- 78
        53121 => X"4F",  -- 79
        53122 => X"50",  -- 80
        53123 => X"50",  -- 80
        53124 => X"50",  -- 80
        53125 => X"51",  -- 81
        53126 => X"53",  -- 83
        53127 => X"55",  -- 85
        53128 => X"56",  -- 86
        53129 => X"53",  -- 83
        53130 => X"4D",  -- 77
        53131 => X"48",  -- 72
        53132 => X"4B",  -- 75
        53133 => X"52",  -- 82
        53134 => X"54",  -- 84
        53135 => X"51",  -- 81
        53136 => X"49",  -- 73
        53137 => X"49",  -- 73
        53138 => X"49",  -- 73
        53139 => X"48",  -- 72
        53140 => X"48",  -- 72
        53141 => X"45",  -- 69
        53142 => X"40",  -- 64
        53143 => X"3D",  -- 61
        53144 => X"3A",  -- 58
        53145 => X"30",  -- 48
        53146 => X"46",  -- 70
        53147 => X"5F",  -- 95
        53148 => X"4E",  -- 78
        53149 => X"34",  -- 52
        53150 => X"2D",  -- 45
        53151 => X"2C",  -- 44
        53152 => X"31",  -- 49
        53153 => X"30",  -- 48
        53154 => X"30",  -- 48
        53155 => X"32",  -- 50
        53156 => X"32",  -- 50
        53157 => X"30",  -- 48
        53158 => X"32",  -- 50
        53159 => X"36",  -- 54
        53160 => X"27",  -- 39
        53161 => X"2F",  -- 47
        53162 => X"40",  -- 64
        53163 => X"39",  -- 57
        53164 => X"30",  -- 48
        53165 => X"36",  -- 54
        53166 => X"40",  -- 64
        53167 => X"53",  -- 83
        53168 => X"5E",  -- 94
        53169 => X"52",  -- 82
        53170 => X"4F",  -- 79
        53171 => X"4F",  -- 79
        53172 => X"4A",  -- 74
        53173 => X"45",  -- 69
        53174 => X"45",  -- 69
        53175 => X"47",  -- 71
        53176 => X"53",  -- 83
        53177 => X"63",  -- 99
        53178 => X"69",  -- 105
        53179 => X"50",  -- 80
        53180 => X"49",  -- 73
        53181 => X"43",  -- 67
        53182 => X"27",  -- 39
        53183 => X"28",  -- 40
        53184 => X"1D",  -- 29
        53185 => X"1F",  -- 31
        53186 => X"4C",  -- 76
        53187 => X"56",  -- 86
        53188 => X"48",  -- 72
        53189 => X"52",  -- 82
        53190 => X"4B",  -- 75
        53191 => X"36",  -- 54
        53192 => X"37",  -- 55
        53193 => X"4B",  -- 75
        53194 => X"43",  -- 67
        53195 => X"31",  -- 49
        53196 => X"38",  -- 56
        53197 => X"42",  -- 66
        53198 => X"3F",  -- 63
        53199 => X"3D",  -- 61
        53200 => X"3D",  -- 61
        53201 => X"4B",  -- 75
        53202 => X"68",  -- 104
        53203 => X"66",  -- 102
        53204 => X"62",  -- 98
        53205 => X"6A",  -- 106
        53206 => X"66",  -- 102
        53207 => X"73",  -- 115
        53208 => X"70",  -- 112
        53209 => X"70",  -- 112
        53210 => X"72",  -- 114
        53211 => X"76",  -- 118
        53212 => X"78",  -- 120
        53213 => X"75",  -- 117
        53214 => X"6F",  -- 111
        53215 => X"69",  -- 105
        53216 => X"70",  -- 112
        53217 => X"6B",  -- 107
        53218 => X"7D",  -- 125
        53219 => X"7D",  -- 125
        53220 => X"77",  -- 119
        53221 => X"80",  -- 128
        53222 => X"7B",  -- 123
        53223 => X"73",  -- 115
        53224 => X"67",  -- 103
        53225 => X"5B",  -- 91
        53226 => X"59",  -- 89
        53227 => X"5E",  -- 94
        53228 => X"83",  -- 131
        53229 => X"75",  -- 117
        53230 => X"63",  -- 99
        53231 => X"69",  -- 105
        53232 => X"66",  -- 102
        53233 => X"60",  -- 96
        53234 => X"63",  -- 99
        53235 => X"72",  -- 114
        53236 => X"80",  -- 128
        53237 => X"82",  -- 130
        53238 => X"7F",  -- 127
        53239 => X"7C",  -- 124
        53240 => X"3D",  -- 61
        53241 => X"5D",  -- 93
        53242 => X"8D",  -- 141
        53243 => X"8C",  -- 140
        53244 => X"6C",  -- 108
        53245 => X"40",  -- 64
        53246 => X"59",  -- 89
        53247 => X"86",  -- 134
        53248 => X"85",  -- 133
        53249 => X"B7",  -- 183
        53250 => X"D3",  -- 211
        53251 => X"9A",  -- 154
        53252 => X"6B",  -- 107
        53253 => X"60",  -- 96
        53254 => X"5A",  -- 90
        53255 => X"5E",  -- 94
        53256 => X"63",  -- 99
        53257 => X"74",  -- 116
        53258 => X"74",  -- 116
        53259 => X"6E",  -- 110
        53260 => X"6C",  -- 108
        53261 => X"62",  -- 98
        53262 => X"5F",  -- 95
        53263 => X"6A",  -- 106
        53264 => X"6D",  -- 109
        53265 => X"72",  -- 114
        53266 => X"6F",  -- 111
        53267 => X"7D",  -- 125
        53268 => X"77",  -- 119
        53269 => X"76",  -- 118
        53270 => X"73",  -- 115
        53271 => X"61",  -- 97
        53272 => X"7E",  -- 126
        53273 => X"A4",  -- 164
        53274 => X"96",  -- 150
        53275 => X"73",  -- 115
        53276 => X"71",  -- 113
        53277 => X"55",  -- 85
        53278 => X"4F",  -- 79
        53279 => X"70",  -- 112
        53280 => X"5D",  -- 93
        53281 => X"85",  -- 133
        53282 => X"88",  -- 136
        53283 => X"8E",  -- 142
        53284 => X"97",  -- 151
        53285 => X"81",  -- 129
        53286 => X"45",  -- 69
        53287 => X"1C",  -- 28
        53288 => X"20",  -- 32
        53289 => X"14",  -- 20
        53290 => X"2A",  -- 42
        53291 => X"37",  -- 55
        53292 => X"33",  -- 51
        53293 => X"2D",  -- 45
        53294 => X"22",  -- 34
        53295 => X"2C",  -- 44
        53296 => X"32",  -- 50
        53297 => X"34",  -- 52
        53298 => X"3A",  -- 58
        53299 => X"3D",  -- 61
        53300 => X"3B",  -- 59
        53301 => X"38",  -- 56
        53302 => X"3A",  -- 58
        53303 => X"40",  -- 64
        53304 => X"43",  -- 67
        53305 => X"40",  -- 64
        53306 => X"3B",  -- 59
        53307 => X"3A",  -- 58
        53308 => X"3B",  -- 59
        53309 => X"3A",  -- 58
        53310 => X"39",  -- 57
        53311 => X"38",  -- 56
        53312 => X"39",  -- 57
        53313 => X"3F",  -- 63
        53314 => X"44",  -- 68
        53315 => X"44",  -- 68
        53316 => X"3F",  -- 63
        53317 => X"3D",  -- 61
        53318 => X"40",  -- 64
        53319 => X"44",  -- 68
        53320 => X"55",  -- 85
        53321 => X"61",  -- 97
        53322 => X"6E",  -- 110
        53323 => X"74",  -- 116
        53324 => X"75",  -- 117
        53325 => X"75",  -- 117
        53326 => X"74",  -- 116
        53327 => X"72",  -- 114
        53328 => X"67",  -- 103
        53329 => X"5A",  -- 90
        53330 => X"4F",  -- 79
        53331 => X"48",  -- 72
        53332 => X"45",  -- 69
        53333 => X"42",  -- 66
        53334 => X"43",  -- 67
        53335 => X"47",  -- 71
        53336 => X"4D",  -- 77
        53337 => X"42",  -- 66
        53338 => X"51",  -- 81
        53339 => X"65",  -- 101
        53340 => X"7D",  -- 125
        53341 => X"86",  -- 134
        53342 => X"83",  -- 131
        53343 => X"8C",  -- 140
        53344 => X"97",  -- 151
        53345 => X"8C",  -- 140
        53346 => X"95",  -- 149
        53347 => X"91",  -- 145
        53348 => X"95",  -- 149
        53349 => X"8E",  -- 142
        53350 => X"9A",  -- 154
        53351 => X"96",  -- 150
        53352 => X"88",  -- 136
        53353 => X"89",  -- 137
        53354 => X"97",  -- 151
        53355 => X"A0",  -- 160
        53356 => X"97",  -- 151
        53357 => X"92",  -- 146
        53358 => X"97",  -- 151
        53359 => X"9A",  -- 154
        53360 => X"93",  -- 147
        53361 => X"9D",  -- 157
        53362 => X"A0",  -- 160
        53363 => X"98",  -- 152
        53364 => X"A4",  -- 164
        53365 => X"A0",  -- 160
        53366 => X"A0",  -- 160
        53367 => X"AA",  -- 170
        53368 => X"AF",  -- 175
        53369 => X"B4",  -- 180
        53370 => X"AD",  -- 173
        53371 => X"9C",  -- 156
        53372 => X"A6",  -- 166
        53373 => X"A0",  -- 160
        53374 => X"A3",  -- 163
        53375 => X"89",  -- 137
        53376 => X"9B",  -- 155
        53377 => X"9F",  -- 159
        53378 => X"93",  -- 147
        53379 => X"9B",  -- 155
        53380 => X"A6",  -- 166
        53381 => X"A5",  -- 165
        53382 => X"AF",  -- 175
        53383 => X"B3",  -- 179
        53384 => X"AB",  -- 171
        53385 => X"BD",  -- 189
        53386 => X"B5",  -- 181
        53387 => X"B1",  -- 177
        53388 => X"C2",  -- 194
        53389 => X"C4",  -- 196
        53390 => X"C0",  -- 192
        53391 => X"CC",  -- 204
        53392 => X"D4",  -- 212
        53393 => X"D3",  -- 211
        53394 => X"C5",  -- 197
        53395 => X"AC",  -- 172
        53396 => X"9D",  -- 157
        53397 => X"9D",  -- 157
        53398 => X"A2",  -- 162
        53399 => X"A2",  -- 162
        53400 => X"AD",  -- 173
        53401 => X"A6",  -- 166
        53402 => X"A4",  -- 164
        53403 => X"A9",  -- 169
        53404 => X"AD",  -- 173
        53405 => X"AC",  -- 172
        53406 => X"AA",  -- 170
        53407 => X"A9",  -- 169
        53408 => X"B2",  -- 178
        53409 => X"A9",  -- 169
        53410 => X"A3",  -- 163
        53411 => X"A5",  -- 165
        53412 => X"A5",  -- 165
        53413 => X"9C",  -- 156
        53414 => X"8E",  -- 142
        53415 => X"85",  -- 133
        53416 => X"82",  -- 130
        53417 => X"77",  -- 119
        53418 => X"65",  -- 101
        53419 => X"60",  -- 96
        53420 => X"6A",  -- 106
        53421 => X"6C",  -- 108
        53422 => X"60",  -- 96
        53423 => X"55",  -- 85
        53424 => X"43",  -- 67
        53425 => X"3E",  -- 62
        53426 => X"40",  -- 64
        53427 => X"48",  -- 72
        53428 => X"4C",  -- 76
        53429 => X"4F",  -- 79
        53430 => X"5B",  -- 91
        53431 => X"6A",  -- 106
        53432 => X"73",  -- 115
        53433 => X"70",  -- 112
        53434 => X"73",  -- 115
        53435 => X"81",  -- 129
        53436 => X"8E",  -- 142
        53437 => X"96",  -- 150
        53438 => X"9A",  -- 154
        53439 => X"9D",  -- 157
        53440 => X"51",  -- 81
        53441 => X"4F",  -- 79
        53442 => X"4C",  -- 76
        53443 => X"49",  -- 73
        53444 => X"47",  -- 71
        53445 => X"47",  -- 71
        53446 => X"49",  -- 73
        53447 => X"4A",  -- 74
        53448 => X"49",  -- 73
        53449 => X"45",  -- 69
        53450 => X"3D",  -- 61
        53451 => X"38",  -- 56
        53452 => X"3E",  -- 62
        53453 => X"4A",  -- 74
        53454 => X"4D",  -- 77
        53455 => X"4B",  -- 75
        53456 => X"40",  -- 64
        53457 => X"41",  -- 65
        53458 => X"42",  -- 66
        53459 => X"44",  -- 68
        53460 => X"45",  -- 69
        53461 => X"43",  -- 67
        53462 => X"3B",  -- 59
        53463 => X"35",  -- 53
        53464 => X"2B",  -- 43
        53465 => X"4D",  -- 77
        53466 => X"55",  -- 85
        53467 => X"3F",  -- 63
        53468 => X"31",  -- 49
        53469 => X"34",  -- 52
        53470 => X"34",  -- 52
        53471 => X"30",  -- 48
        53472 => X"36",  -- 54
        53473 => X"34",  -- 52
        53474 => X"34",  -- 52
        53475 => X"36",  -- 54
        53476 => X"31",  -- 49
        53477 => X"2D",  -- 45
        53478 => X"37",  -- 55
        53479 => X"45",  -- 69
        53480 => X"4B",  -- 75
        53481 => X"48",  -- 72
        53482 => X"57",  -- 87
        53483 => X"5F",  -- 95
        53484 => X"6C",  -- 108
        53485 => X"75",  -- 117
        53486 => X"65",  -- 101
        53487 => X"5F",  -- 95
        53488 => X"56",  -- 86
        53489 => X"4F",  -- 79
        53490 => X"4C",  -- 76
        53491 => X"4B",  -- 75
        53492 => X"53",  -- 83
        53493 => X"6C",  -- 108
        53494 => X"7A",  -- 122
        53495 => X"76",  -- 118
        53496 => X"65",  -- 101
        53497 => X"45",  -- 69
        53498 => X"37",  -- 55
        53499 => X"3C",  -- 60
        53500 => X"51",  -- 81
        53501 => X"50",  -- 80
        53502 => X"3C",  -- 60
        53503 => X"53",  -- 83
        53504 => X"38",  -- 56
        53505 => X"2F",  -- 47
        53506 => X"55",  -- 85
        53507 => X"4D",  -- 77
        53508 => X"2B",  -- 43
        53509 => X"3C",  -- 60
        53510 => X"4C",  -- 76
        53511 => X"46",  -- 70
        53512 => X"52",  -- 82
        53513 => X"5E",  -- 94
        53514 => X"3E",  -- 62
        53515 => X"1D",  -- 29
        53516 => X"2F",  -- 47
        53517 => X"4A",  -- 74
        53518 => X"48",  -- 72
        53519 => X"45",  -- 69
        53520 => X"3F",  -- 63
        53521 => X"44",  -- 68
        53522 => X"5D",  -- 93
        53523 => X"5A",  -- 90
        53524 => X"58",  -- 88
        53525 => X"60",  -- 96
        53526 => X"5E",  -- 94
        53527 => X"6E",  -- 110
        53528 => X"6D",  -- 109
        53529 => X"6E",  -- 110
        53530 => X"6C",  -- 108
        53531 => X"6A",  -- 106
        53532 => X"6F",  -- 111
        53533 => X"76",  -- 118
        53534 => X"77",  -- 119
        53535 => X"75",  -- 117
        53536 => X"72",  -- 114
        53537 => X"63",  -- 99
        53538 => X"79",  -- 121
        53539 => X"81",  -- 129
        53540 => X"6E",  -- 110
        53541 => X"64",  -- 100
        53542 => X"62",  -- 98
        53543 => X"6B",  -- 107
        53544 => X"61",  -- 97
        53545 => X"53",  -- 83
        53546 => X"68",  -- 104
        53547 => X"62",  -- 98
        53548 => X"88",  -- 136
        53549 => X"7B",  -- 123
        53550 => X"52",  -- 82
        53551 => X"60",  -- 96
        53552 => X"7D",  -- 125
        53553 => X"76",  -- 118
        53554 => X"73",  -- 115
        53555 => X"79",  -- 121
        53556 => X"7E",  -- 126
        53557 => X"7B",  -- 123
        53558 => X"75",  -- 117
        53559 => X"72",  -- 114
        53560 => X"3B",  -- 59
        53561 => X"59",  -- 89
        53562 => X"8D",  -- 141
        53563 => X"94",  -- 148
        53564 => X"7C",  -- 124
        53565 => X"5D",  -- 93
        53566 => X"74",  -- 116
        53567 => X"8B",  -- 139
        53568 => X"6E",  -- 110
        53569 => X"B4",  -- 180
        53570 => X"DF",  -- 223
        53571 => X"BC",  -- 188
        53572 => X"81",  -- 129
        53573 => X"81",  -- 129
        53574 => X"74",  -- 116
        53575 => X"88",  -- 136
        53576 => X"75",  -- 117
        53577 => X"8C",  -- 140
        53578 => X"92",  -- 146
        53579 => X"8C",  -- 140
        53580 => X"87",  -- 135
        53581 => X"78",  -- 120
        53582 => X"6F",  -- 111
        53583 => X"7A",  -- 122
        53584 => X"64",  -- 100
        53585 => X"6B",  -- 107
        53586 => X"65",  -- 101
        53587 => X"7D",  -- 125
        53588 => X"7B",  -- 123
        53589 => X"83",  -- 131
        53590 => X"71",  -- 113
        53591 => X"54",  -- 84
        53592 => X"5E",  -- 94
        53593 => X"8A",  -- 138
        53594 => X"76",  -- 118
        53595 => X"7E",  -- 126
        53596 => X"96",  -- 150
        53597 => X"75",  -- 117
        53598 => X"53",  -- 83
        53599 => X"53",  -- 83
        53600 => X"53",  -- 83
        53601 => X"84",  -- 132
        53602 => X"72",  -- 114
        53603 => X"83",  -- 131
        53604 => X"84",  -- 132
        53605 => X"73",  -- 115
        53606 => X"4B",  -- 75
        53607 => X"15",  -- 21
        53608 => X"16",  -- 22
        53609 => X"10",  -- 16
        53610 => X"27",  -- 39
        53611 => X"30",  -- 48
        53612 => X"31",  -- 49
        53613 => X"31",  -- 49
        53614 => X"29",  -- 41
        53615 => X"3B",  -- 59
        53616 => X"33",  -- 51
        53617 => X"36",  -- 54
        53618 => X"39",  -- 57
        53619 => X"3B",  -- 59
        53620 => X"38",  -- 56
        53621 => X"35",  -- 53
        53622 => X"37",  -- 55
        53623 => X"3E",  -- 62
        53624 => X"3A",  -- 58
        53625 => X"37",  -- 55
        53626 => X"34",  -- 52
        53627 => X"35",  -- 53
        53628 => X"3A",  -- 58
        53629 => X"3D",  -- 61
        53630 => X"3B",  -- 59
        53631 => X"38",  -- 56
        53632 => X"3B",  -- 59
        53633 => X"41",  -- 65
        53634 => X"44",  -- 68
        53635 => X"3F",  -- 63
        53636 => X"3A",  -- 58
        53637 => X"3F",  -- 63
        53638 => X"4F",  -- 79
        53639 => X"5F",  -- 95
        53640 => X"6A",  -- 106
        53641 => X"73",  -- 115
        53642 => X"76",  -- 118
        53643 => X"72",  -- 114
        53644 => X"6C",  -- 108
        53645 => X"69",  -- 105
        53646 => X"66",  -- 102
        53647 => X"64",  -- 100
        53648 => X"57",  -- 87
        53649 => X"4C",  -- 76
        53650 => X"44",  -- 68
        53651 => X"46",  -- 70
        53652 => X"48",  -- 72
        53653 => X"46",  -- 70
        53654 => X"44",  -- 68
        53655 => X"45",  -- 69
        53656 => X"44",  -- 68
        53657 => X"41",  -- 65
        53658 => X"5D",  -- 93
        53659 => X"74",  -- 116
        53660 => X"7E",  -- 126
        53661 => X"84",  -- 132
        53662 => X"88",  -- 136
        53663 => X"94",  -- 148
        53664 => X"9B",  -- 155
        53665 => X"8E",  -- 142
        53666 => X"9A",  -- 154
        53667 => X"9E",  -- 158
        53668 => X"A2",  -- 162
        53669 => X"93",  -- 147
        53670 => X"97",  -- 151
        53671 => X"92",  -- 146
        53672 => X"88",  -- 136
        53673 => X"8F",  -- 143
        53674 => X"9E",  -- 158
        53675 => X"A4",  -- 164
        53676 => X"97",  -- 151
        53677 => X"8F",  -- 143
        53678 => X"91",  -- 145
        53679 => X"8F",  -- 143
        53680 => X"8A",  -- 138
        53681 => X"96",  -- 150
        53682 => X"95",  -- 149
        53683 => X"7E",  -- 126
        53684 => X"93",  -- 147
        53685 => X"93",  -- 147
        53686 => X"9A",  -- 154
        53687 => X"9A",  -- 154
        53688 => X"AD",  -- 173
        53689 => X"B5",  -- 181
        53690 => X"AD",  -- 173
        53691 => X"96",  -- 150
        53692 => X"9F",  -- 159
        53693 => X"9E",  -- 158
        53694 => X"AF",  -- 175
        53695 => X"9D",  -- 157
        53696 => X"9F",  -- 159
        53697 => X"A1",  -- 161
        53698 => X"96",  -- 150
        53699 => X"A4",  -- 164
        53700 => X"B2",  -- 178
        53701 => X"AC",  -- 172
        53702 => X"B1",  -- 177
        53703 => X"B6",  -- 182
        53704 => X"B0",  -- 176
        53705 => X"C2",  -- 194
        53706 => X"B9",  -- 185
        53707 => X"B2",  -- 178
        53708 => X"C3",  -- 195
        53709 => X"C3",  -- 195
        53710 => X"BD",  -- 189
        53711 => X"C9",  -- 201
        53712 => X"D6",  -- 214
        53713 => X"D3",  -- 211
        53714 => X"C0",  -- 192
        53715 => X"A6",  -- 166
        53716 => X"99",  -- 153
        53717 => X"9C",  -- 156
        53718 => X"A2",  -- 162
        53719 => X"A0",  -- 160
        53720 => X"AD",  -- 173
        53721 => X"A6",  -- 166
        53722 => X"A2",  -- 162
        53723 => X"A7",  -- 167
        53724 => X"AB",  -- 171
        53725 => X"A8",  -- 168
        53726 => X"A5",  -- 165
        53727 => X"A3",  -- 163
        53728 => X"AB",  -- 171
        53729 => X"A2",  -- 162
        53730 => X"9F",  -- 159
        53731 => X"A5",  -- 165
        53732 => X"A6",  -- 166
        53733 => X"99",  -- 153
        53734 => X"85",  -- 133
        53735 => X"78",  -- 120
        53736 => X"8C",  -- 140
        53737 => X"81",  -- 129
        53738 => X"63",  -- 99
        53739 => X"4F",  -- 79
        53740 => X"5A",  -- 90
        53741 => X"66",  -- 102
        53742 => X"60",  -- 96
        53743 => X"56",  -- 86
        53744 => X"4A",  -- 74
        53745 => X"3F",  -- 63
        53746 => X"35",  -- 53
        53747 => X"39",  -- 57
        53748 => X"4B",  -- 75
        53749 => X"5F",  -- 95
        53750 => X"69",  -- 105
        53751 => X"6B",  -- 107
        53752 => X"78",  -- 120
        53753 => X"6D",  -- 109
        53754 => X"65",  -- 101
        53755 => X"6C",  -- 108
        53756 => X"79",  -- 121
        53757 => X"88",  -- 136
        53758 => X"97",  -- 151
        53759 => X"A2",  -- 162
        53760 => X"46",  -- 70
        53761 => X"44",  -- 68
        53762 => X"41",  -- 65
        53763 => X"3D",  -- 61
        53764 => X"3A",  -- 58
        53765 => X"38",  -- 56
        53766 => X"36",  -- 54
        53767 => X"36",  -- 54
        53768 => X"3E",  -- 62
        53769 => X"38",  -- 56
        53770 => X"33",  -- 51
        53771 => X"31",  -- 49
        53772 => X"33",  -- 51
        53773 => X"36",  -- 54
        53774 => X"38",  -- 56
        53775 => X"37",  -- 55
        53776 => X"36",  -- 54
        53777 => X"31",  -- 49
        53778 => X"2E",  -- 46
        53779 => X"30",  -- 48
        53780 => X"36",  -- 54
        53781 => X"39",  -- 57
        53782 => X"30",  -- 48
        53783 => X"26",  -- 38
        53784 => X"49",  -- 73
        53785 => X"42",  -- 66
        53786 => X"38",  -- 56
        53787 => X"30",  -- 48
        53788 => X"30",  -- 48
        53789 => X"37",  -- 55
        53790 => X"38",  -- 56
        53791 => X"36",  -- 54
        53792 => X"37",  -- 55
        53793 => X"42",  -- 66
        53794 => X"4C",  -- 76
        53795 => X"52",  -- 82
        53796 => X"55",  -- 85
        53797 => X"57",  -- 87
        53798 => X"55",  -- 85
        53799 => X"50",  -- 80
        53800 => X"3A",  -- 58
        53801 => X"39",  -- 57
        53802 => X"38",  -- 56
        53803 => X"32",  -- 50
        53804 => X"26",  -- 38
        53805 => X"22",  -- 34
        53806 => X"26",  -- 38
        53807 => X"26",  -- 38
        53808 => X"21",  -- 33
        53809 => X"1E",  -- 30
        53810 => X"27",  -- 39
        53811 => X"41",  -- 65
        53812 => X"55",  -- 85
        53813 => X"55",  -- 85
        53814 => X"43",  -- 67
        53815 => X"35",  -- 53
        53816 => X"38",  -- 56
        53817 => X"67",  -- 103
        53818 => X"59",  -- 89
        53819 => X"41",  -- 65
        53820 => X"45",  -- 69
        53821 => X"49",  -- 73
        53822 => X"4D",  -- 77
        53823 => X"53",  -- 83
        53824 => X"48",  -- 72
        53825 => X"47",  -- 71
        53826 => X"4C",  -- 76
        53827 => X"4B",  -- 75
        53828 => X"3E",  -- 62
        53829 => X"3A",  -- 58
        53830 => X"45",  -- 69
        53831 => X"4E",  -- 78
        53832 => X"5F",  -- 95
        53833 => X"6D",  -- 109
        53834 => X"43",  -- 67
        53835 => X"15",  -- 21
        53836 => X"27",  -- 39
        53837 => X"45",  -- 69
        53838 => X"48",  -- 72
        53839 => X"4C",  -- 76
        53840 => X"4E",  -- 78
        53841 => X"54",  -- 84
        53842 => X"5C",  -- 92
        53843 => X"62",  -- 98
        53844 => X"5B",  -- 91
        53845 => X"57",  -- 87
        53846 => X"63",  -- 99
        53847 => X"76",  -- 118
        53848 => X"62",  -- 98
        53849 => X"80",  -- 128
        53850 => X"6F",  -- 111
        53851 => X"70",  -- 112
        53852 => X"78",  -- 120
        53853 => X"7A",  -- 122
        53854 => X"69",  -- 105
        53855 => X"87",  -- 135
        53856 => X"64",  -- 100
        53857 => X"66",  -- 102
        53858 => X"6A",  -- 106
        53859 => X"70",  -- 112
        53860 => X"73",  -- 115
        53861 => X"6E",  -- 110
        53862 => X"6A",  -- 106
        53863 => X"66",  -- 102
        53864 => X"69",  -- 105
        53865 => X"67",  -- 103
        53866 => X"66",  -- 102
        53867 => X"64",  -- 100
        53868 => X"7F",  -- 127
        53869 => X"77",  -- 119
        53870 => X"25",  -- 37
        53871 => X"59",  -- 89
        53872 => X"87",  -- 135
        53873 => X"7D",  -- 125
        53874 => X"72",  -- 114
        53875 => X"6E",  -- 110
        53876 => X"7B",  -- 123
        53877 => X"7A",  -- 122
        53878 => X"72",  -- 114
        53879 => X"87",  -- 135
        53880 => X"6C",  -- 108
        53881 => X"95",  -- 149
        53882 => X"9E",  -- 158
        53883 => X"A0",  -- 160
        53884 => X"90",  -- 144
        53885 => X"64",  -- 100
        53886 => X"3F",  -- 63
        53887 => X"89",  -- 137
        53888 => X"BD",  -- 189
        53889 => X"D3",  -- 211
        53890 => X"F0",  -- 240
        53891 => X"DE",  -- 222
        53892 => X"CB",  -- 203
        53893 => X"B9",  -- 185
        53894 => X"BC",  -- 188
        53895 => X"B0",  -- 176
        53896 => X"A1",  -- 161
        53897 => X"9C",  -- 156
        53898 => X"9C",  -- 156
        53899 => X"A3",  -- 163
        53900 => X"9A",  -- 154
        53901 => X"A7",  -- 167
        53902 => X"A5",  -- 165
        53903 => X"BA",  -- 186
        53904 => X"A3",  -- 163
        53905 => X"81",  -- 129
        53906 => X"8B",  -- 139
        53907 => X"7C",  -- 124
        53908 => X"5A",  -- 90
        53909 => X"81",  -- 129
        53910 => X"68",  -- 104
        53911 => X"4A",  -- 74
        53912 => X"5E",  -- 94
        53913 => X"79",  -- 121
        53914 => X"6D",  -- 109
        53915 => X"64",  -- 100
        53916 => X"6F",  -- 111
        53917 => X"97",  -- 151
        53918 => X"7C",  -- 124
        53919 => X"52",  -- 82
        53920 => X"59",  -- 89
        53921 => X"67",  -- 103
        53922 => X"5F",  -- 95
        53923 => X"5B",  -- 91
        53924 => X"6F",  -- 111
        53925 => X"6A",  -- 106
        53926 => X"3B",  -- 59
        53927 => X"13",  -- 19
        53928 => X"0F",  -- 15
        53929 => X"17",  -- 23
        53930 => X"20",  -- 32
        53931 => X"2B",  -- 43
        53932 => X"32",  -- 50
        53933 => X"36",  -- 54
        53934 => X"39",  -- 57
        53935 => X"3B",  -- 59
        53936 => X"3C",  -- 60
        53937 => X"3A",  -- 58
        53938 => X"39",  -- 57
        53939 => X"36",  -- 54
        53940 => X"35",  -- 53
        53941 => X"38",  -- 56
        53942 => X"3A",  -- 58
        53943 => X"3E",  -- 62
        53944 => X"38",  -- 56
        53945 => X"35",  -- 53
        53946 => X"35",  -- 53
        53947 => X"38",  -- 56
        53948 => X"38",  -- 56
        53949 => X"35",  -- 53
        53950 => X"38",  -- 56
        53951 => X"3F",  -- 63
        53952 => X"3C",  -- 60
        53953 => X"43",  -- 67
        53954 => X"45",  -- 69
        53955 => X"3D",  -- 61
        53956 => X"3A",  -- 58
        53957 => X"48",  -- 72
        53958 => X"63",  -- 99
        53959 => X"75",  -- 117
        53960 => X"7C",  -- 124
        53961 => X"77",  -- 119
        53962 => X"74",  -- 116
        53963 => X"72",  -- 114
        53964 => X"6C",  -- 108
        53965 => X"5F",  -- 95
        53966 => X"55",  -- 85
        53967 => X"50",  -- 80
        53968 => X"46",  -- 70
        53969 => X"48",  -- 72
        53970 => X"4A",  -- 74
        53971 => X"49",  -- 73
        53972 => X"46",  -- 70
        53973 => X"44",  -- 68
        53974 => X"44",  -- 68
        53975 => X"45",  -- 69
        53976 => X"40",  -- 64
        53977 => X"41",  -- 65
        53978 => X"59",  -- 89
        53979 => X"79",  -- 121
        53980 => X"88",  -- 136
        53981 => X"8D",  -- 141
        53982 => X"98",  -- 152
        53983 => X"9E",  -- 158
        53984 => X"A4",  -- 164
        53985 => X"A1",  -- 161
        53986 => X"A3",  -- 163
        53987 => X"A8",  -- 168
        53988 => X"A6",  -- 166
        53989 => X"9B",  -- 155
        53990 => X"95",  -- 149
        53991 => X"95",  -- 149
        53992 => X"8C",  -- 140
        53993 => X"A0",  -- 160
        53994 => X"9B",  -- 155
        53995 => X"9A",  -- 154
        53996 => X"9E",  -- 158
        53997 => X"91",  -- 145
        53998 => X"8F",  -- 143
        53999 => X"95",  -- 149
        54000 => X"8D",  -- 141
        54001 => X"9E",  -- 158
        54002 => X"99",  -- 153
        54003 => X"8A",  -- 138
        54004 => X"8F",  -- 143
        54005 => X"95",  -- 149
        54006 => X"9C",  -- 156
        54007 => X"AA",  -- 170
        54008 => X"AC",  -- 172
        54009 => X"B7",  -- 183
        54010 => X"B0",  -- 176
        54011 => X"A6",  -- 166
        54012 => X"A9",  -- 169
        54013 => X"9F",  -- 159
        54014 => X"95",  -- 149
        54015 => X"9A",  -- 154
        54016 => X"B6",  -- 182
        54017 => X"AE",  -- 174
        54018 => X"A9",  -- 169
        54019 => X"AE",  -- 174
        54020 => X"B4",  -- 180
        54021 => X"B4",  -- 180
        54022 => X"B3",  -- 179
        54023 => X"B7",  -- 183
        54024 => X"B6",  -- 182
        54025 => X"B6",  -- 182
        54026 => X"B8",  -- 184
        54027 => X"BE",  -- 190
        54028 => X"C4",  -- 196
        54029 => X"C9",  -- 201
        54030 => X"C9",  -- 201
        54031 => X"C8",  -- 200
        54032 => X"CC",  -- 204
        54033 => X"CD",  -- 205
        54034 => X"B5",  -- 181
        54035 => X"94",  -- 148
        54036 => X"A0",  -- 160
        54037 => X"94",  -- 148
        54038 => X"A2",  -- 162
        54039 => X"A2",  -- 162
        54040 => X"A9",  -- 169
        54041 => X"A7",  -- 167
        54042 => X"A8",  -- 168
        54043 => X"A7",  -- 167
        54044 => X"A5",  -- 165
        54045 => X"A7",  -- 167
        54046 => X"A2",  -- 162
        54047 => X"90",  -- 144
        54048 => X"99",  -- 153
        54049 => X"AC",  -- 172
        54050 => X"A4",  -- 164
        54051 => X"96",  -- 150
        54052 => X"92",  -- 146
        54053 => X"9F",  -- 159
        54054 => X"97",  -- 151
        54055 => X"68",  -- 104
        54056 => X"6B",  -- 107
        54057 => X"8B",  -- 139
        54058 => X"7A",  -- 122
        54059 => X"5B",  -- 91
        54060 => X"45",  -- 69
        54061 => X"49",  -- 73
        54062 => X"62",  -- 98
        54063 => X"55",  -- 85
        54064 => X"45",  -- 69
        54065 => X"48",  -- 72
        54066 => X"45",  -- 69
        54067 => X"45",  -- 69
        54068 => X"4E",  -- 78
        54069 => X"5F",  -- 95
        54070 => X"6B",  -- 107
        54071 => X"6F",  -- 111
        54072 => X"71",  -- 113
        54073 => X"7E",  -- 126
        54074 => X"77",  -- 119
        54075 => X"64",  -- 100
        54076 => X"61",  -- 97
        54077 => X"6E",  -- 110
        54078 => X"81",  -- 129
        54079 => X"92",  -- 146
        54080 => X"3A",  -- 58
        54081 => X"39",  -- 57
        54082 => X"37",  -- 55
        54083 => X"36",  -- 54
        54084 => X"33",  -- 51
        54085 => X"32",  -- 50
        54086 => X"31",  -- 49
        54087 => X"30",  -- 48
        54088 => X"34",  -- 52
        54089 => X"33",  -- 51
        54090 => X"31",  -- 49
        54091 => X"2F",  -- 47
        54092 => X"2A",  -- 42
        54093 => X"2A",  -- 42
        54094 => X"2D",  -- 45
        54095 => X"2F",  -- 47
        54096 => X"2C",  -- 44
        54097 => X"2D",  -- 45
        54098 => X"2E",  -- 46
        54099 => X"2B",  -- 43
        54100 => X"2A",  -- 42
        54101 => X"2D",  -- 45
        54102 => X"36",  -- 54
        54103 => X"3E",  -- 62
        54104 => X"39",  -- 57
        54105 => X"33",  -- 51
        54106 => X"2E",  -- 46
        54107 => X"31",  -- 49
        54108 => X"2F",  -- 47
        54109 => X"2D",  -- 45
        54110 => X"30",  -- 48
        54111 => X"36",  -- 54
        54112 => X"42",  -- 66
        54113 => X"46",  -- 70
        54114 => X"47",  -- 71
        54115 => X"3F",  -- 63
        54116 => X"37",  -- 55
        54117 => X"32",  -- 50
        54118 => X"2A",  -- 42
        54119 => X"22",  -- 34
        54120 => X"39",  -- 57
        54121 => X"2B",  -- 43
        54122 => X"24",  -- 36
        54123 => X"25",  -- 37
        54124 => X"23",  -- 35
        54125 => X"23",  -- 35
        54126 => X"20",  -- 32
        54127 => X"18",  -- 24
        54128 => X"29",  -- 41
        54129 => X"49",  -- 73
        54130 => X"58",  -- 88
        54131 => X"43",  -- 67
        54132 => X"27",  -- 39
        54133 => X"23",  -- 35
        54134 => X"31",  -- 49
        54135 => X"3B",  -- 59
        54136 => X"2B",  -- 43
        54137 => X"87",  -- 135
        54138 => X"7D",  -- 125
        54139 => X"42",  -- 66
        54140 => X"3B",  -- 59
        54141 => X"3B",  -- 59
        54142 => X"3E",  -- 62
        54143 => X"52",  -- 82
        54144 => X"54",  -- 84
        54145 => X"53",  -- 83
        54146 => X"51",  -- 81
        54147 => X"4D",  -- 77
        54148 => X"46",  -- 70
        54149 => X"4C",  -- 76
        54150 => X"57",  -- 87
        54151 => X"5D",  -- 93
        54152 => X"66",  -- 102
        54153 => X"6D",  -- 109
        54154 => X"50",  -- 80
        54155 => X"1F",  -- 31
        54156 => X"1A",  -- 26
        54157 => X"3F",  -- 63
        54158 => X"57",  -- 87
        54159 => X"54",  -- 84
        54160 => X"43",  -- 67
        54161 => X"50",  -- 80
        54162 => X"61",  -- 97
        54163 => X"69",  -- 105
        54164 => X"65",  -- 101
        54165 => X"61",  -- 97
        54166 => X"67",  -- 103
        54167 => X"71",  -- 113
        54168 => X"65",  -- 101
        54169 => X"7B",  -- 123
        54170 => X"7C",  -- 124
        54171 => X"67",  -- 103
        54172 => X"66",  -- 102
        54173 => X"6B",  -- 107
        54174 => X"6F",  -- 111
        54175 => X"6D",  -- 109
        54176 => X"7F",  -- 127
        54177 => X"79",  -- 121
        54178 => X"76",  -- 118
        54179 => X"76",  -- 118
        54180 => X"77",  -- 119
        54181 => X"78",  -- 120
        54182 => X"7F",  -- 127
        54183 => X"87",  -- 135
        54184 => X"88",  -- 136
        54185 => X"7A",  -- 122
        54186 => X"85",  -- 133
        54187 => X"83",  -- 131
        54188 => X"78",  -- 120
        54189 => X"59",  -- 89
        54190 => X"0F",  -- 15
        54191 => X"2A",  -- 42
        54192 => X"7E",  -- 126
        54193 => X"89",  -- 137
        54194 => X"7F",  -- 127
        54195 => X"68",  -- 104
        54196 => X"67",  -- 103
        54197 => X"6F",  -- 111
        54198 => X"74",  -- 116
        54199 => X"82",  -- 130
        54200 => X"98",  -- 152
        54201 => X"8E",  -- 142
        54202 => X"9F",  -- 159
        54203 => X"9E",  -- 158
        54204 => X"92",  -- 146
        54205 => X"68",  -- 104
        54206 => X"3B",  -- 59
        54207 => X"7A",  -- 122
        54208 => X"AA",  -- 170
        54209 => X"C9",  -- 201
        54210 => X"E0",  -- 224
        54211 => X"C1",  -- 193
        54212 => X"9F",  -- 159
        54213 => X"74",  -- 116
        54214 => X"67",  -- 103
        54215 => X"5A",  -- 90
        54216 => X"67",  -- 103
        54217 => X"62",  -- 98
        54218 => X"63",  -- 99
        54219 => X"6A",  -- 106
        54220 => X"5F",  -- 95
        54221 => X"66",  -- 102
        54222 => X"5A",  -- 90
        54223 => X"68",  -- 104
        54224 => X"68",  -- 104
        54225 => X"74",  -- 116
        54226 => X"9D",  -- 157
        54227 => X"B1",  -- 177
        54228 => X"9D",  -- 157
        54229 => X"9A",  -- 154
        54230 => X"77",  -- 119
        54231 => X"45",  -- 69
        54232 => X"42",  -- 66
        54233 => X"75",  -- 117
        54234 => X"76",  -- 118
        54235 => X"72",  -- 114
        54236 => X"7D",  -- 125
        54237 => X"6B",  -- 107
        54238 => X"5D",  -- 93
        54239 => X"8A",  -- 138
        54240 => X"68",  -- 104
        54241 => X"6B",  -- 107
        54242 => X"5E",  -- 94
        54243 => X"56",  -- 86
        54244 => X"5C",  -- 92
        54245 => X"50",  -- 80
        54246 => X"36",  -- 54
        54247 => X"26",  -- 38
        54248 => X"16",  -- 22
        54249 => X"19",  -- 25
        54250 => X"1E",  -- 30
        54251 => X"28",  -- 40
        54252 => X"33",  -- 51
        54253 => X"3A",  -- 58
        54254 => X"3F",  -- 63
        54255 => X"41",  -- 65
        54256 => X"40",  -- 64
        54257 => X"3D",  -- 61
        54258 => X"3A",  -- 58
        54259 => X"36",  -- 54
        54260 => X"36",  -- 54
        54261 => X"39",  -- 57
        54262 => X"40",  -- 64
        54263 => X"44",  -- 68
        54264 => X"3C",  -- 60
        54265 => X"37",  -- 55
        54266 => X"35",  -- 53
        54267 => X"38",  -- 56
        54268 => X"37",  -- 55
        54269 => X"37",  -- 55
        54270 => X"38",  -- 56
        54271 => X"3D",  -- 61
        54272 => X"3E",  -- 62
        54273 => X"43",  -- 67
        54274 => X"44",  -- 68
        54275 => X"3F",  -- 63
        54276 => X"41",  -- 65
        54277 => X"52",  -- 82
        54278 => X"6A",  -- 106
        54279 => X"7C",  -- 124
        54280 => X"83",  -- 131
        54281 => X"7A",  -- 122
        54282 => X"71",  -- 113
        54283 => X"6E",  -- 110
        54284 => X"69",  -- 105
        54285 => X"5E",  -- 94
        54286 => X"54",  -- 84
        54287 => X"4F",  -- 79
        54288 => X"45",  -- 69
        54289 => X"48",  -- 72
        54290 => X"4C",  -- 76
        54291 => X"4D",  -- 77
        54292 => X"4B",  -- 75
        54293 => X"49",  -- 73
        54294 => X"45",  -- 69
        54295 => X"45",  -- 69
        54296 => X"40",  -- 64
        54297 => X"4F",  -- 79
        54298 => X"62",  -- 98
        54299 => X"74",  -- 116
        54300 => X"86",  -- 134
        54301 => X"93",  -- 147
        54302 => X"9C",  -- 156
        54303 => X"9F",  -- 159
        54304 => X"A3",  -- 163
        54305 => X"A6",  -- 166
        54306 => X"A9",  -- 169
        54307 => X"AB",  -- 171
        54308 => X"AB",  -- 171
        54309 => X"A3",  -- 163
        54310 => X"94",  -- 148
        54311 => X"86",  -- 134
        54312 => X"92",  -- 146
        54313 => X"98",  -- 152
        54314 => X"93",  -- 147
        54315 => X"8F",  -- 143
        54316 => X"9C",  -- 156
        54317 => X"9E",  -- 158
        54318 => X"92",  -- 146
        54319 => X"94",  -- 148
        54320 => X"88",  -- 136
        54321 => X"93",  -- 147
        54322 => X"96",  -- 150
        54323 => X"90",  -- 144
        54324 => X"8E",  -- 142
        54325 => X"8C",  -- 140
        54326 => X"8D",  -- 141
        54327 => X"96",  -- 150
        54328 => X"A4",  -- 164
        54329 => X"AA",  -- 170
        54330 => X"A5",  -- 165
        54331 => X"9E",  -- 158
        54332 => X"A0",  -- 160
        54333 => X"9E",  -- 158
        54334 => X"98",  -- 152
        54335 => X"96",  -- 150
        54336 => X"A8",  -- 168
        54337 => X"AC",  -- 172
        54338 => X"AF",  -- 175
        54339 => X"B0",  -- 176
        54340 => X"B1",  -- 177
        54341 => X"B3",  -- 179
        54342 => X"B5",  -- 181
        54343 => X"B8",  -- 184
        54344 => X"BF",  -- 191
        54345 => X"BE",  -- 190
        54346 => X"BE",  -- 190
        54347 => X"C0",  -- 192
        54348 => X"C2",  -- 194
        54349 => X"C6",  -- 198
        54350 => X"C7",  -- 199
        54351 => X"C9",  -- 201
        54352 => X"CD",  -- 205
        54353 => X"CB",  -- 203
        54354 => X"AF",  -- 175
        54355 => X"92",  -- 146
        54356 => X"9D",  -- 157
        54357 => X"91",  -- 145
        54358 => X"9E",  -- 158
        54359 => X"9F",  -- 159
        54360 => X"A7",  -- 167
        54361 => X"A7",  -- 167
        54362 => X"A5",  -- 165
        54363 => X"9E",  -- 158
        54364 => X"A1",  -- 161
        54365 => X"AD",  -- 173
        54366 => X"A6",  -- 166
        54367 => X"8B",  -- 139
        54368 => X"88",  -- 136
        54369 => X"98",  -- 152
        54370 => X"9A",  -- 154
        54371 => X"94",  -- 148
        54372 => X"86",  -- 134
        54373 => X"85",  -- 133
        54374 => X"8F",  -- 143
        54375 => X"81",  -- 129
        54376 => X"5B",  -- 91
        54377 => X"60",  -- 96
        54378 => X"71",  -- 113
        54379 => X"6F",  -- 111
        54380 => X"56",  -- 86
        54381 => X"3E",  -- 62
        54382 => X"3F",  -- 63
        54383 => X"56",  -- 86
        54384 => X"45",  -- 69
        54385 => X"48",  -- 72
        54386 => X"4A",  -- 74
        54387 => X"4D",  -- 77
        54388 => X"56",  -- 86
        54389 => X"65",  -- 101
        54390 => X"6F",  -- 111
        54391 => X"72",  -- 114
        54392 => X"7A",  -- 122
        54393 => X"82",  -- 130
        54394 => X"7F",  -- 127
        54395 => X"73",  -- 115
        54396 => X"6B",  -- 107
        54397 => X"66",  -- 102
        54398 => X"6D",  -- 109
        54399 => X"7F",  -- 127
        54400 => X"36",  -- 54
        54401 => X"36",  -- 54
        54402 => X"36",  -- 54
        54403 => X"35",  -- 53
        54404 => X"35",  -- 53
        54405 => X"33",  -- 51
        54406 => X"32",  -- 50
        54407 => X"32",  -- 50
        54408 => X"2F",  -- 47
        54409 => X"34",  -- 52
        54410 => X"38",  -- 56
        54411 => X"35",  -- 53
        54412 => X"2C",  -- 44
        54413 => X"28",  -- 40
        54414 => X"2B",  -- 43
        54415 => X"30",  -- 48
        54416 => X"2A",  -- 42
        54417 => X"2B",  -- 43
        54418 => X"2F",  -- 47
        54419 => X"31",  -- 49
        54420 => X"2C",  -- 44
        54421 => X"2B",  -- 43
        54422 => X"37",  -- 55
        54423 => X"47",  -- 71
        54424 => X"31",  -- 49
        54425 => X"28",  -- 40
        54426 => X"25",  -- 37
        54427 => X"2A",  -- 42
        54428 => X"27",  -- 39
        54429 => X"21",  -- 33
        54430 => X"28",  -- 40
        54431 => X"39",  -- 57
        54432 => X"40",  -- 64
        54433 => X"42",  -- 66
        54434 => X"42",  -- 66
        54435 => X"3E",  -- 62
        54436 => X"39",  -- 57
        54437 => X"36",  -- 54
        54438 => X"34",  -- 52
        54439 => X"32",  -- 50
        54440 => X"2C",  -- 44
        54441 => X"2E",  -- 46
        54442 => X"21",  -- 33
        54443 => X"26",  -- 38
        54444 => X"30",  -- 48
        54445 => X"1B",  -- 27
        54446 => X"1B",  -- 27
        54447 => X"44",  -- 68
        54448 => X"5F",  -- 95
        54449 => X"47",  -- 71
        54450 => X"28",  -- 40
        54451 => X"18",  -- 24
        54452 => X"27",  -- 39
        54453 => X"3D",  -- 61
        54454 => X"39",  -- 57
        54455 => X"24",  -- 36
        54456 => X"49",  -- 73
        54457 => X"84",  -- 132
        54458 => X"96",  -- 150
        54459 => X"5F",  -- 95
        54460 => X"1E",  -- 30
        54461 => X"23",  -- 35
        54462 => X"4D",  -- 77
        54463 => X"48",  -- 72
        54464 => X"47",  -- 71
        54465 => X"53",  -- 83
        54466 => X"5B",  -- 91
        54467 => X"52",  -- 82
        54468 => X"4A",  -- 74
        54469 => X"4F",  -- 79
        54470 => X"5A",  -- 90
        54471 => X"60",  -- 96
        54472 => X"6D",  -- 109
        54473 => X"89",  -- 137
        54474 => X"7D",  -- 125
        54475 => X"37",  -- 55
        54476 => X"09",  -- 9
        54477 => X"2F",  -- 47
        54478 => X"57",  -- 87
        54479 => X"4B",  -- 75
        54480 => X"5E",  -- 94
        54481 => X"5E",  -- 94
        54482 => X"5B",  -- 91
        54483 => X"57",  -- 87
        54484 => X"5A",  -- 90
        54485 => X"65",  -- 101
        54486 => X"71",  -- 113
        54487 => X"76",  -- 118
        54488 => X"71",  -- 113
        54489 => X"72",  -- 114
        54490 => X"81",  -- 129
        54491 => X"69",  -- 105
        54492 => X"65",  -- 101
        54493 => X"68",  -- 104
        54494 => X"81",  -- 129
        54495 => X"73",  -- 115
        54496 => X"76",  -- 118
        54497 => X"71",  -- 113
        54498 => X"6F",  -- 111
        54499 => X"76",  -- 118
        54500 => X"78",  -- 120
        54501 => X"79",  -- 121
        54502 => X"86",  -- 134
        54503 => X"97",  -- 151
        54504 => X"88",  -- 136
        54505 => X"8F",  -- 143
        54506 => X"8D",  -- 141
        54507 => X"81",  -- 129
        54508 => X"73",  -- 115
        54509 => X"3A",  -- 58
        54510 => X"05",  -- 5
        54511 => X"57",  -- 87
        54512 => X"A3",  -- 163
        54513 => X"A4",  -- 164
        54514 => X"8F",  -- 143
        54515 => X"73",  -- 115
        54516 => X"6E",  -- 110
        54517 => X"76",  -- 118
        54518 => X"80",  -- 128
        54519 => X"88",  -- 136
        54520 => X"95",  -- 149
        54521 => X"8E",  -- 142
        54522 => X"97",  -- 151
        54523 => X"66",  -- 102
        54524 => X"76",  -- 118
        54525 => X"9F",  -- 159
        54526 => X"96",  -- 150
        54527 => X"B2",  -- 178
        54528 => X"C4",  -- 196
        54529 => X"D5",  -- 213
        54530 => X"D3",  -- 211
        54531 => X"AC",  -- 172
        54532 => X"9F",  -- 159
        54533 => X"88",  -- 136
        54534 => X"88",  -- 136
        54535 => X"8D",  -- 141
        54536 => X"8D",  -- 141
        54537 => X"89",  -- 137
        54538 => X"8D",  -- 141
        54539 => X"96",  -- 150
        54540 => X"8C",  -- 140
        54541 => X"92",  -- 146
        54542 => X"85",  -- 133
        54543 => X"92",  -- 146
        54544 => X"7F",  -- 127
        54545 => X"7B",  -- 123
        54546 => X"70",  -- 112
        54547 => X"66",  -- 102
        54548 => X"65",  -- 101
        54549 => X"72",  -- 114
        54550 => X"96",  -- 150
        54551 => X"93",  -- 147
        54552 => X"61",  -- 97
        54553 => X"6D",  -- 109
        54554 => X"6E",  -- 110
        54555 => X"71",  -- 113
        54556 => X"84",  -- 132
        54557 => X"69",  -- 105
        54558 => X"4E",  -- 78
        54559 => X"51",  -- 81
        54560 => X"6D",  -- 109
        54561 => X"76",  -- 118
        54562 => X"6A",  -- 106
        54563 => X"55",  -- 85
        54564 => X"52",  -- 82
        54565 => X"4B",  -- 75
        54566 => X"2D",  -- 45
        54567 => X"12",  -- 18
        54568 => X"1E",  -- 30
        54569 => X"1E",  -- 30
        54570 => X"1E",  -- 30
        54571 => X"26",  -- 38
        54572 => X"2F",  -- 47
        54573 => X"3A",  -- 58
        54574 => X"41",  -- 65
        54575 => X"44",  -- 68
        54576 => X"44",  -- 68
        54577 => X"41",  -- 65
        54578 => X"3C",  -- 60
        54579 => X"39",  -- 57
        54580 => X"39",  -- 57
        54581 => X"3F",  -- 63
        54582 => X"47",  -- 71
        54583 => X"4D",  -- 77
        54584 => X"44",  -- 68
        54585 => X"3F",  -- 63
        54586 => X"3B",  -- 59
        54587 => X"3C",  -- 60
        54588 => X"3C",  -- 60
        54589 => X"3D",  -- 61
        54590 => X"3F",  -- 63
        54591 => X"42",  -- 66
        54592 => X"46",  -- 70
        54593 => X"48",  -- 72
        54594 => X"46",  -- 70
        54595 => X"42",  -- 66
        54596 => X"46",  -- 70
        54597 => X"59",  -- 89
        54598 => X"71",  -- 113
        54599 => X"80",  -- 128
        54600 => X"88",  -- 136
        54601 => X"7C",  -- 124
        54602 => X"72",  -- 114
        54603 => X"6E",  -- 110
        54604 => X"69",  -- 105
        54605 => X"5E",  -- 94
        54606 => X"51",  -- 81
        54607 => X"48",  -- 72
        54608 => X"43",  -- 67
        54609 => X"45",  -- 69
        54610 => X"4B",  -- 75
        54611 => X"4D",  -- 77
        54612 => X"4A",  -- 74
        54613 => X"47",  -- 71
        54614 => X"42",  -- 66
        54615 => X"3F",  -- 63
        54616 => X"3D",  -- 61
        54617 => X"5F",  -- 95
        54618 => X"6F",  -- 111
        54619 => X"73",  -- 115
        54620 => X"88",  -- 136
        54621 => X"9D",  -- 157
        54622 => X"A3",  -- 163
        54623 => X"A6",  -- 166
        54624 => X"A4",  -- 164
        54625 => X"AC",  -- 172
        54626 => X"AE",  -- 174
        54627 => X"AC",  -- 172
        54628 => X"AB",  -- 171
        54629 => X"A6",  -- 166
        54630 => X"92",  -- 146
        54631 => X"7D",  -- 125
        54632 => X"94",  -- 148
        54633 => X"93",  -- 147
        54634 => X"97",  -- 151
        54635 => X"89",  -- 137
        54636 => X"94",  -- 148
        54637 => X"A3",  -- 163
        54638 => X"92",  -- 146
        54639 => X"95",  -- 149
        54640 => X"8E",  -- 142
        54641 => X"8A",  -- 138
        54642 => X"93",  -- 147
        54643 => X"9C",  -- 156
        54644 => X"99",  -- 153
        54645 => X"97",  -- 151
        54646 => X"94",  -- 148
        54647 => X"8F",  -- 143
        54648 => X"8F",  -- 143
        54649 => X"99",  -- 153
        54650 => X"A4",  -- 164
        54651 => X"A0",  -- 160
        54652 => X"94",  -- 148
        54653 => X"95",  -- 149
        54654 => X"98",  -- 152
        54655 => X"92",  -- 146
        54656 => X"9D",  -- 157
        54657 => X"A5",  -- 165
        54658 => X"A8",  -- 168
        54659 => X"A7",  -- 167
        54660 => X"A7",  -- 167
        54661 => X"B0",  -- 176
        54662 => X"BB",  -- 187
        54663 => X"C1",  -- 193
        54664 => X"C2",  -- 194
        54665 => X"C3",  -- 195
        54666 => X"C3",  -- 195
        54667 => X"C1",  -- 193
        54668 => X"C0",  -- 192
        54669 => X"C3",  -- 195
        54670 => X"C7",  -- 199
        54671 => X"CB",  -- 203
        54672 => X"CD",  -- 205
        54673 => X"C7",  -- 199
        54674 => X"A6",  -- 166
        54675 => X"8F",  -- 143
        54676 => X"97",  -- 151
        54677 => X"8E",  -- 142
        54678 => X"97",  -- 151
        54679 => X"9C",  -- 156
        54680 => X"9F",  -- 159
        54681 => X"A7",  -- 167
        54682 => X"A6",  -- 166
        54683 => X"98",  -- 152
        54684 => X"98",  -- 152
        54685 => X"AA",  -- 170
        54686 => X"A8",  -- 168
        54687 => X"8E",  -- 142
        54688 => X"7A",  -- 122
        54689 => X"84",  -- 132
        54690 => X"8F",  -- 143
        54691 => X"96",  -- 150
        54692 => X"7D",  -- 125
        54693 => X"6A",  -- 106
        54694 => X"7E",  -- 126
        54695 => X"8D",  -- 141
        54696 => X"68",  -- 104
        54697 => X"42",  -- 66
        54698 => X"51",  -- 81
        54699 => X"61",  -- 97
        54700 => X"62",  -- 98
        54701 => X"4C",  -- 76
        54702 => X"2D",  -- 45
        54703 => X"43",  -- 67
        54704 => X"4A",  -- 74
        54705 => X"4E",  -- 78
        54706 => X"54",  -- 84
        54707 => X"56",  -- 86
        54708 => X"5C",  -- 92
        54709 => X"66",  -- 102
        54710 => X"6C",  -- 108
        54711 => X"6F",  -- 111
        54712 => X"74",  -- 116
        54713 => X"78",  -- 120
        54714 => X"7A",  -- 122
        54715 => X"7B",  -- 123
        54716 => X"75",  -- 117
        54717 => X"65",  -- 101
        54718 => X"64",  -- 100
        54719 => X"76",  -- 118
        54720 => X"3B",  -- 59
        54721 => X"3A",  -- 58
        54722 => X"3B",  -- 59
        54723 => X"3A",  -- 58
        54724 => X"39",  -- 57
        54725 => X"37",  -- 55
        54726 => X"35",  -- 53
        54727 => X"34",  -- 52
        54728 => X"2E",  -- 46
        54729 => X"35",  -- 53
        54730 => X"3B",  -- 59
        54731 => X"3C",  -- 60
        54732 => X"37",  -- 55
        54733 => X"30",  -- 48
        54734 => X"2E",  -- 46
        54735 => X"2F",  -- 47
        54736 => X"2F",  -- 47
        54737 => X"2F",  -- 47
        54738 => X"37",  -- 55
        54739 => X"41",  -- 65
        54740 => X"3E",  -- 62
        54741 => X"31",  -- 49
        54742 => X"2D",  -- 45
        54743 => X"32",  -- 50
        54744 => X"2F",  -- 47
        54745 => X"2B",  -- 43
        54746 => X"26",  -- 38
        54747 => X"23",  -- 35
        54748 => X"1F",  -- 31
        54749 => X"1F",  -- 31
        54750 => X"2D",  -- 45
        54751 => X"3E",  -- 62
        54752 => X"41",  -- 65
        54753 => X"40",  -- 64
        54754 => X"3B",  -- 59
        54755 => X"36",  -- 54
        54756 => X"32",  -- 50
        54757 => X"31",  -- 49
        54758 => X"31",  -- 49
        54759 => X"33",  -- 51
        54760 => X"27",  -- 39
        54761 => X"2A",  -- 42
        54762 => X"2C",  -- 44
        54763 => X"2A",  -- 42
        54764 => X"24",  -- 36
        54765 => X"27",  -- 39
        54766 => X"3F",  -- 63
        54767 => X"5E",  -- 94
        54768 => X"3E",  -- 62
        54769 => X"2F",  -- 47
        54770 => X"27",  -- 39
        54771 => X"27",  -- 39
        54772 => X"27",  -- 39
        54773 => X"28",  -- 40
        54774 => X"32",  -- 50
        54775 => X"3E",  -- 62
        54776 => X"2D",  -- 45
        54777 => X"61",  -- 97
        54778 => X"A1",  -- 161
        54779 => X"8D",  -- 141
        54780 => X"3E",  -- 62
        54781 => X"4A",  -- 74
        54782 => X"6B",  -- 107
        54783 => X"2E",  -- 46
        54784 => X"1C",  -- 28
        54785 => X"40",  -- 64
        54786 => X"56",  -- 86
        54787 => X"51",  -- 81
        54788 => X"49",  -- 73
        54789 => X"4D",  -- 77
        54790 => X"59",  -- 89
        54791 => X"62",  -- 98
        54792 => X"7A",  -- 122
        54793 => X"9B",  -- 155
        54794 => X"A1",  -- 161
        54795 => X"65",  -- 101
        54796 => X"22",  -- 34
        54797 => X"15",  -- 21
        54798 => X"31",  -- 49
        54799 => X"47",  -- 71
        54800 => X"55",  -- 85
        54801 => X"54",  -- 84
        54802 => X"53",  -- 83
        54803 => X"53",  -- 83
        54804 => X"60",  -- 96
        54805 => X"6B",  -- 107
        54806 => X"69",  -- 105
        54807 => X"5F",  -- 95
        54808 => X"68",  -- 104
        54809 => X"64",  -- 100
        54810 => X"7C",  -- 124
        54811 => X"85",  -- 133
        54812 => X"85",  -- 133
        54813 => X"75",  -- 117
        54814 => X"79",  -- 121
        54815 => X"73",  -- 115
        54816 => X"6D",  -- 109
        54817 => X"71",  -- 113
        54818 => X"7A",  -- 122
        54819 => X"87",  -- 135
        54820 => X"86",  -- 134
        54821 => X"80",  -- 128
        54822 => X"83",  -- 131
        54823 => X"90",  -- 144
        54824 => X"81",  -- 129
        54825 => X"85",  -- 133
        54826 => X"7F",  -- 127
        54827 => X"6A",  -- 106
        54828 => X"49",  -- 73
        54829 => X"14",  -- 20
        54830 => X"1C",  -- 28
        54831 => X"93",  -- 147
        54832 => X"C2",  -- 194
        54833 => X"B2",  -- 178
        54834 => X"95",  -- 149
        54835 => X"8B",  -- 139
        54836 => X"83",  -- 131
        54837 => X"7D",  -- 125
        54838 => X"89",  -- 137
        54839 => X"95",  -- 149
        54840 => X"8E",  -- 142
        54841 => X"9A",  -- 154
        54842 => X"7B",  -- 123
        54843 => X"2C",  -- 44
        54844 => X"66",  -- 102
        54845 => X"BF",  -- 191
        54846 => X"CA",  -- 202
        54847 => X"B1",  -- 177
        54848 => X"B8",  -- 184
        54849 => X"D2",  -- 210
        54850 => X"D3",  -- 211
        54851 => X"B0",  -- 176
        54852 => X"A6",  -- 166
        54853 => X"87",  -- 135
        54854 => X"7E",  -- 126
        54855 => X"86",  -- 134
        54856 => X"7F",  -- 127
        54857 => X"7D",  -- 125
        54858 => X"83",  -- 131
        54859 => X"8C",  -- 140
        54860 => X"82",  -- 130
        54861 => X"89",  -- 137
        54862 => X"80",  -- 128
        54863 => X"92",  -- 146
        54864 => X"92",  -- 146
        54865 => X"A0",  -- 160
        54866 => X"AE",  -- 174
        54867 => X"A3",  -- 163
        54868 => X"9D",  -- 157
        54869 => X"7C",  -- 124
        54870 => X"6D",  -- 109
        54871 => X"5E",  -- 94
        54872 => X"8C",  -- 140
        54873 => X"9C",  -- 156
        54874 => X"7B",  -- 123
        54875 => X"5B",  -- 91
        54876 => X"7E",  -- 126
        54877 => X"5A",  -- 90
        54878 => X"3A",  -- 58
        54879 => X"54",  -- 84
        54880 => X"45",  -- 69
        54881 => X"60",  -- 96
        54882 => X"6E",  -- 110
        54883 => X"60",  -- 96
        54884 => X"4C",  -- 76
        54885 => X"3E",  -- 62
        54886 => X"32",  -- 50
        54887 => X"2C",  -- 44
        54888 => X"22",  -- 34
        54889 => X"22",  -- 34
        54890 => X"21",  -- 33
        54891 => X"24",  -- 36
        54892 => X"2A",  -- 42
        54893 => X"33",  -- 51
        54894 => X"3A",  -- 58
        54895 => X"40",  -- 64
        54896 => X"42",  -- 66
        54897 => X"40",  -- 64
        54898 => X"3D",  -- 61
        54899 => X"3B",  -- 59
        54900 => X"3D",  -- 61
        54901 => X"44",  -- 68
        54902 => X"4E",  -- 78
        54903 => X"54",  -- 84
        54904 => X"4E",  -- 78
        54905 => X"49",  -- 73
        54906 => X"45",  -- 69
        54907 => X"45",  -- 69
        54908 => X"47",  -- 71
        54909 => X"4A",  -- 74
        54910 => X"4C",  -- 76
        54911 => X"4C",  -- 76
        54912 => X"4E",  -- 78
        54913 => X"4D",  -- 77
        54914 => X"49",  -- 73
        54915 => X"44",  -- 68
        54916 => X"4B",  -- 75
        54917 => X"5F",  -- 95
        54918 => X"71",  -- 113
        54919 => X"7C",  -- 124
        54920 => X"83",  -- 131
        54921 => X"7E",  -- 126
        54922 => X"7A",  -- 122
        54923 => X"76",  -- 118
        54924 => X"6C",  -- 108
        54925 => X"5B",  -- 91
        54926 => X"4A",  -- 74
        54927 => X"42",  -- 66
        54928 => X"44",  -- 68
        54929 => X"47",  -- 71
        54930 => X"4A",  -- 74
        54931 => X"4B",  -- 75
        54932 => X"47",  -- 71
        54933 => X"42",  -- 66
        54934 => X"40",  -- 64
        54935 => X"3D",  -- 61
        54936 => X"3F",  -- 63
        54937 => X"6B",  -- 107
        54938 => X"7A",  -- 122
        54939 => X"7F",  -- 127
        54940 => X"99",  -- 153
        54941 => X"AA",  -- 170
        54942 => X"AC",  -- 172
        54943 => X"B6",  -- 182
        54944 => X"B0",  -- 176
        54945 => X"B1",  -- 177
        54946 => X"B0",  -- 176
        54947 => X"AF",  -- 175
        54948 => X"AC",  -- 172
        54949 => X"A5",  -- 165
        54950 => X"95",  -- 149
        54951 => X"89",  -- 137
        54952 => X"90",  -- 144
        54953 => X"90",  -- 144
        54954 => X"A4",  -- 164
        54955 => X"90",  -- 144
        54956 => X"8E",  -- 142
        54957 => X"A4",  -- 164
        54958 => X"94",  -- 148
        54959 => X"9F",  -- 159
        54960 => X"A1",  -- 161
        54961 => X"8D",  -- 141
        54962 => X"8F",  -- 143
        54963 => X"9D",  -- 157
        54964 => X"9E",  -- 158
        54965 => X"9E",  -- 158
        54966 => X"9B",  -- 155
        54967 => X"90",  -- 144
        54968 => X"8A",  -- 138
        54969 => X"8B",  -- 139
        54970 => X"95",  -- 149
        54971 => X"97",  -- 151
        54972 => X"8D",  -- 141
        54973 => X"8E",  -- 142
        54974 => X"89",  -- 137
        54975 => X"72",  -- 114
        54976 => X"84",  -- 132
        54977 => X"87",  -- 135
        54978 => X"8F",  -- 143
        54979 => X"9A",  -- 154
        54980 => X"A6",  -- 166
        54981 => X"B0",  -- 176
        54982 => X"BC",  -- 188
        54983 => X"C4",  -- 196
        54984 => X"BE",  -- 190
        54985 => X"C1",  -- 193
        54986 => X"C4",  -- 196
        54987 => X"C3",  -- 195
        54988 => X"C1",  -- 193
        54989 => X"C2",  -- 194
        54990 => X"C7",  -- 199
        54991 => X"CD",  -- 205
        54992 => X"CD",  -- 205
        54993 => X"C3",  -- 195
        54994 => X"9D",  -- 157
        54995 => X"8C",  -- 140
        54996 => X"95",  -- 149
        54997 => X"8C",  -- 140
        54998 => X"91",  -- 145
        54999 => X"99",  -- 153
        55000 => X"96",  -- 150
        55001 => X"A3",  -- 163
        55002 => X"A7",  -- 167
        55003 => X"99",  -- 153
        55004 => X"8F",  -- 143
        55005 => X"9A",  -- 154
        55006 => X"A2",  -- 162
        55007 => X"97",  -- 151
        55008 => X"79",  -- 121
        55009 => X"79",  -- 121
        55010 => X"80",  -- 128
        55011 => X"8D",  -- 141
        55012 => X"75",  -- 117
        55013 => X"59",  -- 89
        55014 => X"65",  -- 101
        55015 => X"72",  -- 114
        55016 => X"79",  -- 121
        55017 => X"50",  -- 80
        55018 => X"3B",  -- 59
        55019 => X"3C",  -- 60
        55020 => X"50",  -- 80
        55021 => X"57",  -- 87
        55022 => X"3F",  -- 63
        55023 => X"38",  -- 56
        55024 => X"47",  -- 71
        55025 => X"4C",  -- 76
        55026 => X"53",  -- 83
        55027 => X"58",  -- 88
        55028 => X"5C",  -- 92
        55029 => X"63",  -- 99
        55030 => X"6B",  -- 107
        55031 => X"70",  -- 112
        55032 => X"6D",  -- 109
        55033 => X"6F",  -- 111
        55034 => X"6E",  -- 110
        55035 => X"71",  -- 113
        55036 => X"71",  -- 113
        55037 => X"66",  -- 102
        55038 => X"62",  -- 98
        55039 => X"6D",  -- 109
        55040 => X"38",  -- 56
        55041 => X"38",  -- 56
        55042 => X"39",  -- 57
        55043 => X"38",  -- 56
        55044 => X"36",  -- 54
        55045 => X"33",  -- 51
        55046 => X"30",  -- 48
        55047 => X"2F",  -- 47
        55048 => X"2D",  -- 45
        55049 => X"2F",  -- 47
        55050 => X"35",  -- 53
        55051 => X"38",  -- 56
        55052 => X"37",  -- 55
        55053 => X"32",  -- 50
        55054 => X"28",  -- 40
        55055 => X"21",  -- 33
        55056 => X"2A",  -- 42
        55057 => X"34",  -- 52
        55058 => X"42",  -- 66
        55059 => X"4B",  -- 75
        55060 => X"40",  -- 64
        55061 => X"2B",  -- 43
        55062 => X"1F",  -- 31
        55063 => X"1D",  -- 29
        55064 => X"2D",  -- 45
        55065 => X"31",  -- 49
        55066 => X"2F",  -- 47
        55067 => X"26",  -- 38
        55068 => X"23",  -- 35
        55069 => X"2D",  -- 45
        55070 => X"39",  -- 57
        55071 => X"3D",  -- 61
        55072 => X"36",  -- 54
        55073 => X"33",  -- 51
        55074 => X"2C",  -- 44
        55075 => X"28",  -- 40
        55076 => X"24",  -- 36
        55077 => X"25",  -- 37
        55078 => X"29",  -- 41
        55079 => X"2D",  -- 45
        55080 => X"2E",  -- 46
        55081 => X"1A",  -- 26
        55082 => X"22",  -- 34
        55083 => X"1D",  -- 29
        55084 => X"14",  -- 20
        55085 => X"44",  -- 68
        55086 => X"5F",  -- 95
        55087 => X"33",  -- 51
        55088 => X"34",  -- 52
        55089 => X"28",  -- 40
        55090 => X"25",  -- 37
        55091 => X"31",  -- 49
        55092 => X"37",  -- 55
        55093 => X"2E",  -- 46
        55094 => X"26",  -- 38
        55095 => X"22",  -- 34
        55096 => X"1A",  -- 26
        55097 => X"68",  -- 104
        55098 => X"9C",  -- 156
        55099 => X"86",  -- 134
        55100 => X"5C",  -- 92
        55101 => X"66",  -- 102
        55102 => X"6C",  -- 108
        55103 => X"2D",  -- 45
        55104 => X"0B",  -- 11
        55105 => X"2A",  -- 42
        55106 => X"3A",  -- 58
        55107 => X"39",  -- 57
        55108 => X"41",  -- 65
        55109 => X"50",  -- 80
        55110 => X"61",  -- 97
        55111 => X"74",  -- 116
        55112 => X"8A",  -- 138
        55113 => X"9A",  -- 154
        55114 => X"A0",  -- 160
        55115 => X"92",  -- 146
        55116 => X"5F",  -- 95
        55117 => X"16",  -- 22
        55118 => X"0B",  -- 11
        55119 => X"41",  -- 65
        55120 => X"3A",  -- 58
        55121 => X"41",  -- 65
        55122 => X"45",  -- 69
        55123 => X"48",  -- 72
        55124 => X"53",  -- 83
        55125 => X"5F",  -- 95
        55126 => X"63",  -- 99
        55127 => X"60",  -- 96
        55128 => X"75",  -- 117
        55129 => X"74",  -- 116
        55130 => X"6E",  -- 110
        55131 => X"7C",  -- 124
        55132 => X"7E",  -- 126
        55133 => X"7A",  -- 122
        55134 => X"6D",  -- 109
        55135 => X"7C",  -- 124
        55136 => X"78",  -- 120
        55137 => X"7E",  -- 126
        55138 => X"85",  -- 133
        55139 => X"89",  -- 137
        55140 => X"7E",  -- 126
        55141 => X"6F",  -- 111
        55142 => X"6B",  -- 107
        55143 => X"70",  -- 112
        55144 => X"68",  -- 104
        55145 => X"4A",  -- 74
        55146 => X"59",  -- 89
        55147 => X"48",  -- 72
        55148 => X"0B",  -- 11
        55149 => X"14",  -- 20
        55150 => X"71",  -- 113
        55151 => X"B1",  -- 177
        55152 => X"BC",  -- 188
        55153 => X"AF",  -- 175
        55154 => X"96",  -- 150
        55155 => X"94",  -- 148
        55156 => X"88",  -- 136
        55157 => X"78",  -- 120
        55158 => X"81",  -- 129
        55159 => X"81",  -- 129
        55160 => X"85",  -- 133
        55161 => X"9A",  -- 154
        55162 => X"66",  -- 102
        55163 => X"4D",  -- 77
        55164 => X"9F",  -- 159
        55165 => X"C8",  -- 200
        55166 => X"C7",  -- 199
        55167 => X"98",  -- 152
        55168 => X"78",  -- 120
        55169 => X"9B",  -- 155
        55170 => X"A7",  -- 167
        55171 => X"88",  -- 136
        55172 => X"7C",  -- 124
        55173 => X"5A",  -- 90
        55174 => X"55",  -- 85
        55175 => X"64",  -- 100
        55176 => X"5A",  -- 90
        55177 => X"5D",  -- 93
        55178 => X"67",  -- 103
        55179 => X"6F",  -- 111
        55180 => X"5F",  -- 95
        55181 => X"61",  -- 97
        55182 => X"59",  -- 89
        55183 => X"6B",  -- 107
        55184 => X"51",  -- 81
        55185 => X"4D",  -- 77
        55186 => X"61",  -- 97
        55187 => X"4E",  -- 78
        55188 => X"66",  -- 102
        55189 => X"75",  -- 117
        55190 => X"78",  -- 120
        55191 => X"8E",  -- 142
        55192 => X"8C",  -- 140
        55193 => X"7D",  -- 125
        55194 => X"A6",  -- 166
        55195 => X"B7",  -- 183
        55196 => X"97",  -- 151
        55197 => X"5E",  -- 94
        55198 => X"4D",  -- 77
        55199 => X"38",  -- 56
        55200 => X"3C",  -- 60
        55201 => X"41",  -- 65
        55202 => X"56",  -- 86
        55203 => X"6B",  -- 107
        55204 => X"66",  -- 102
        55205 => X"49",  -- 73
        55206 => X"29",  -- 41
        55207 => X"15",  -- 21
        55208 => X"1B",  -- 27
        55209 => X"1F",  -- 31
        55210 => X"22",  -- 34
        55211 => X"24",  -- 36
        55212 => X"27",  -- 39
        55213 => X"2C",  -- 44
        55214 => X"33",  -- 51
        55215 => X"39",  -- 57
        55216 => X"3B",  -- 59
        55217 => X"3B",  -- 59
        55218 => X"3C",  -- 60
        55219 => X"3D",  -- 61
        55220 => X"40",  -- 64
        55221 => X"47",  -- 71
        55222 => X"50",  -- 80
        55223 => X"55",  -- 85
        55224 => X"53",  -- 83
        55225 => X"4F",  -- 79
        55226 => X"4B",  -- 75
        55227 => X"4C",  -- 76
        55228 => X"51",  -- 81
        55229 => X"57",  -- 87
        55230 => X"58",  -- 88
        55231 => X"55",  -- 85
        55232 => X"52",  -- 82
        55233 => X"51",  -- 81
        55234 => X"4D",  -- 77
        55235 => X"4A",  -- 74
        55236 => X"53",  -- 83
        55237 => X"63",  -- 99
        55238 => X"72",  -- 114
        55239 => X"7A",  -- 122
        55240 => X"7F",  -- 127
        55241 => X"7E",  -- 126
        55242 => X"7B",  -- 123
        55243 => X"75",  -- 117
        55244 => X"66",  -- 102
        55245 => X"54",  -- 84
        55246 => X"46",  -- 70
        55247 => X"43",  -- 67
        55248 => X"48",  -- 72
        55249 => X"49",  -- 73
        55250 => X"49",  -- 73
        55251 => X"48",  -- 72
        55252 => X"43",  -- 67
        55253 => X"40",  -- 64
        55254 => X"40",  -- 64
        55255 => X"3F",  -- 63
        55256 => X"4C",  -- 76
        55257 => X"74",  -- 116
        55258 => X"87",  -- 135
        55259 => X"95",  -- 149
        55260 => X"AD",  -- 173
        55261 => X"B2",  -- 178
        55262 => X"B0",  -- 176
        55263 => X"BE",  -- 190
        55264 => X"B7",  -- 183
        55265 => X"B3",  -- 179
        55266 => X"B6",  -- 182
        55267 => X"BB",  -- 187
        55268 => X"B4",  -- 180
        55269 => X"A3",  -- 163
        55270 => X"99",  -- 153
        55271 => X"9B",  -- 155
        55272 => X"89",  -- 137
        55273 => X"87",  -- 135
        55274 => X"A5",  -- 165
        55275 => X"96",  -- 150
        55276 => X"97",  -- 151
        55277 => X"AD",  -- 173
        55278 => X"9D",  -- 157
        55279 => X"A4",  -- 164
        55280 => X"AD",  -- 173
        55281 => X"98",  -- 152
        55282 => X"96",  -- 150
        55283 => X"97",  -- 151
        55284 => X"8F",  -- 143
        55285 => X"8E",  -- 142
        55286 => X"95",  -- 149
        55287 => X"93",  -- 147
        55288 => X"AA",  -- 170
        55289 => X"97",  -- 151
        55290 => X"92",  -- 146
        55291 => X"98",  -- 152
        55292 => X"9C",  -- 156
        55293 => X"A3",  -- 163
        55294 => X"94",  -- 148
        55295 => X"74",  -- 116
        55296 => X"73",  -- 115
        55297 => X"6F",  -- 111
        55298 => X"7B",  -- 123
        55299 => X"98",  -- 152
        55300 => X"AD",  -- 173
        55301 => X"B2",  -- 178
        55302 => X"B6",  -- 182
        55303 => X"BC",  -- 188
        55304 => X"BB",  -- 187
        55305 => X"C0",  -- 192
        55306 => X"C6",  -- 198
        55307 => X"C6",  -- 198
        55308 => X"C3",  -- 195
        55309 => X"C3",  -- 195
        55310 => X"C6",  -- 198
        55311 => X"CD",  -- 205
        55312 => X"CE",  -- 206
        55313 => X"BF",  -- 191
        55314 => X"93",  -- 147
        55315 => X"8C",  -- 140
        55316 => X"91",  -- 145
        55317 => X"89",  -- 137
        55318 => X"8A",  -- 138
        55319 => X"95",  -- 149
        55320 => X"9A",  -- 154
        55321 => X"99",  -- 153
        55322 => X"9C",  -- 156
        55323 => X"97",  -- 151
        55324 => X"8D",  -- 141
        55325 => X"90",  -- 144
        55326 => X"99",  -- 153
        55327 => X"96",  -- 150
        55328 => X"83",  -- 131
        55329 => X"76",  -- 118
        55330 => X"6D",  -- 109
        55331 => X"74",  -- 116
        55332 => X"66",  -- 102
        55333 => X"52",  -- 82
        55334 => X"53",  -- 83
        55335 => X"4C",  -- 76
        55336 => X"67",  -- 103
        55337 => X"63",  -- 99
        55338 => X"44",  -- 68
        55339 => X"34",  -- 52
        55340 => X"37",  -- 55
        55341 => X"44",  -- 68
        55342 => X"53",  -- 83
        55343 => X"46",  -- 70
        55344 => X"3C",  -- 60
        55345 => X"41",  -- 65
        55346 => X"4A",  -- 74
        55347 => X"50",  -- 80
        55348 => X"57",  -- 87
        55349 => X"60",  -- 96
        55350 => X"6E",  -- 110
        55351 => X"79",  -- 121
        55352 => X"76",  -- 118
        55353 => X"75",  -- 117
        55354 => X"69",  -- 105
        55355 => X"5E",  -- 94
        55356 => X"5F",  -- 95
        55357 => X"5B",  -- 91
        55358 => X"56",  -- 86
        55359 => X"59",  -- 89
        55360 => X"34",  -- 52
        55361 => X"34",  -- 52
        55362 => X"33",  -- 51
        55363 => X"30",  -- 48
        55364 => X"30",  -- 48
        55365 => X"2D",  -- 45
        55366 => X"2C",  -- 44
        55367 => X"2A",  -- 42
        55368 => X"2D",  -- 45
        55369 => X"2B",  -- 43
        55370 => X"2B",  -- 43
        55371 => X"2F",  -- 47
        55372 => X"32",  -- 50
        55373 => X"2E",  -- 46
        55374 => X"21",  -- 33
        55375 => X"15",  -- 21
        55376 => X"20",  -- 32
        55377 => X"35",  -- 53
        55378 => X"48",  -- 72
        55379 => X"47",  -- 71
        55380 => X"32",  -- 50
        55381 => X"20",  -- 32
        55382 => X"1A",  -- 26
        55383 => X"1C",  -- 28
        55384 => X"25",  -- 37
        55385 => X"31",  -- 49
        55386 => X"34",  -- 52
        55387 => X"2E",  -- 46
        55388 => X"2F",  -- 47
        55389 => X"3A",  -- 58
        55390 => X"3B",  -- 59
        55391 => X"34",  -- 52
        55392 => X"27",  -- 39
        55393 => X"24",  -- 36
        55394 => X"21",  -- 33
        55395 => X"20",  -- 32
        55396 => X"22",  -- 34
        55397 => X"26",  -- 38
        55398 => X"2E",  -- 46
        55399 => X"37",  -- 55
        55400 => X"2D",  -- 45
        55401 => X"23",  -- 35
        55402 => X"0F",  -- 15
        55403 => X"15",  -- 21
        55404 => X"35",  -- 53
        55405 => X"3C",  -- 60
        55406 => X"30",  -- 48
        55407 => X"2E",  -- 46
        55408 => X"3B",  -- 59
        55409 => X"3E",  -- 62
        55410 => X"3A",  -- 58
        55411 => X"2C",  -- 44
        55412 => X"23",  -- 35
        55413 => X"24",  -- 36
        55414 => X"26",  -- 38
        55415 => X"26",  -- 38
        55416 => X"2D",  -- 45
        55417 => X"48",  -- 72
        55418 => X"74",  -- 116
        55419 => X"80",  -- 128
        55420 => X"55",  -- 85
        55421 => X"54",  -- 84
        55422 => X"70",  -- 112
        55423 => X"5A",  -- 90
        55424 => X"2C",  -- 44
        55425 => X"34",  -- 52
        55426 => X"25",  -- 37
        55427 => X"1A",  -- 26
        55428 => X"2C",  -- 44
        55429 => X"43",  -- 67
        55430 => X"58",  -- 88
        55431 => X"71",  -- 113
        55432 => X"8B",  -- 139
        55433 => X"A6",  -- 166
        55434 => X"A4",  -- 164
        55435 => X"97",  -- 151
        55436 => X"82",  -- 130
        55437 => X"46",  -- 70
        55438 => X"17",  -- 23
        55439 => X"1E",  -- 30
        55440 => X"2B",  -- 43
        55441 => X"36",  -- 54
        55442 => X"3F",  -- 63
        55443 => X"3D",  -- 61
        55444 => X"3E",  -- 62
        55445 => X"49",  -- 73
        55446 => X"5D",  -- 93
        55447 => X"6C",  -- 108
        55448 => X"77",  -- 119
        55449 => X"81",  -- 129
        55450 => X"6B",  -- 107
        55451 => X"6D",  -- 109
        55452 => X"6D",  -- 109
        55453 => X"7F",  -- 127
        55454 => X"77",  -- 119
        55455 => X"86",  -- 134
        55456 => X"76",  -- 118
        55457 => X"7A",  -- 122
        55458 => X"79",  -- 121
        55459 => X"6C",  -- 108
        55460 => X"5D",  -- 93
        55461 => X"54",  -- 84
        55462 => X"51",  -- 81
        55463 => X"50",  -- 80
        55464 => X"4B",  -- 75
        55465 => X"34",  -- 52
        55466 => X"2B",  -- 43
        55467 => X"13",  -- 19
        55468 => X"0C",  -- 12
        55469 => X"4A",  -- 74
        55470 => X"B4",  -- 180
        55471 => X"CB",  -- 203
        55472 => X"C6",  -- 198
        55473 => X"B7",  -- 183
        55474 => X"94",  -- 148
        55475 => X"8D",  -- 141
        55476 => X"86",  -- 134
        55477 => X"7A",  -- 122
        55478 => X"70",  -- 112
        55479 => X"43",  -- 67
        55480 => X"55",  -- 85
        55481 => X"93",  -- 147
        55482 => X"83",  -- 131
        55483 => X"8F",  -- 143
        55484 => X"B9",  -- 185
        55485 => X"BB",  -- 187
        55486 => X"D2",  -- 210
        55487 => X"BA",  -- 186
        55488 => X"95",  -- 149
        55489 => X"95",  -- 149
        55490 => X"85",  -- 133
        55491 => X"62",  -- 98
        55492 => X"62",  -- 98
        55493 => X"59",  -- 89
        55494 => X"64",  -- 100
        55495 => X"70",  -- 112
        55496 => X"4C",  -- 76
        55497 => X"54",  -- 84
        55498 => X"64",  -- 100
        55499 => X"71",  -- 113
        55500 => X"61",  -- 97
        55501 => X"5E",  -- 94
        55502 => X"4E",  -- 78
        55503 => X"5A",  -- 90
        55504 => X"50",  -- 80
        55505 => X"4B",  -- 75
        55506 => X"62",  -- 98
        55507 => X"48",  -- 72
        55508 => X"4D",  -- 77
        55509 => X"53",  -- 83
        55510 => X"34",  -- 52
        55511 => X"39",  -- 57
        55512 => X"45",  -- 69
        55513 => X"5F",  -- 95
        55514 => X"87",  -- 135
        55515 => X"A1",  -- 161
        55516 => X"AB",  -- 171
        55517 => X"8E",  -- 142
        55518 => X"70",  -- 112
        55519 => X"61",  -- 97
        55520 => X"46",  -- 70
        55521 => X"41",  -- 65
        55522 => X"42",  -- 66
        55523 => X"4A",  -- 74
        55524 => X"58",  -- 88
        55525 => X"65",  -- 101
        55526 => X"50",  -- 80
        55527 => X"27",  -- 39
        55528 => X"17",  -- 23
        55529 => X"1B",  -- 27
        55530 => X"1F",  -- 31
        55531 => X"24",  -- 36
        55532 => X"28",  -- 40
        55533 => X"2D",  -- 45
        55534 => X"34",  -- 52
        55535 => X"39",  -- 57
        55536 => X"35",  -- 53
        55537 => X"37",  -- 55
        55538 => X"3A",  -- 58
        55539 => X"3D",  -- 61
        55540 => X"3F",  -- 63
        55541 => X"45",  -- 69
        55542 => X"4C",  -- 76
        55543 => X"51",  -- 81
        55544 => X"52",  -- 82
        55545 => X"4F",  -- 79
        55546 => X"4C",  -- 76
        55547 => X"4E",  -- 78
        55548 => X"56",  -- 86
        55549 => X"5D",  -- 93
        55550 => X"5D",  -- 93
        55551 => X"57",  -- 87
        55552 => X"50",  -- 80
        55553 => X"51",  -- 81
        55554 => X"4F",  -- 79
        55555 => X"4F",  -- 79
        55556 => X"58",  -- 88
        55557 => X"65",  -- 101
        55558 => X"70",  -- 112
        55559 => X"76",  -- 118
        55560 => X"78",  -- 120
        55561 => X"76",  -- 118
        55562 => X"72",  -- 114
        55563 => X"67",  -- 103
        55564 => X"58",  -- 88
        55565 => X"49",  -- 73
        55566 => X"46",  -- 70
        55567 => X"4B",  -- 75
        55568 => X"49",  -- 73
        55569 => X"47",  -- 71
        55570 => X"46",  -- 70
        55571 => X"42",  -- 66
        55572 => X"3F",  -- 63
        55573 => X"3D",  -- 61
        55574 => X"3D",  -- 61
        55575 => X"40",  -- 64
        55576 => X"5C",  -- 92
        55577 => X"78",  -- 120
        55578 => X"8F",  -- 143
        55579 => X"A3",  -- 163
        55580 => X"B3",  -- 179
        55581 => X"AD",  -- 173
        55582 => X"A6",  -- 166
        55583 => X"B1",  -- 177
        55584 => X"AF",  -- 175
        55585 => X"AA",  -- 170
        55586 => X"B1",  -- 177
        55587 => X"BD",  -- 189
        55588 => X"B5",  -- 181
        55589 => X"9E",  -- 158
        55590 => X"95",  -- 149
        55591 => X"9C",  -- 156
        55592 => X"8A",  -- 138
        55593 => X"81",  -- 129
        55594 => X"96",  -- 150
        55595 => X"9A",  -- 154
        55596 => X"A4",  -- 164
        55597 => X"B4",  -- 180
        55598 => X"A7",  -- 167
        55599 => X"9F",  -- 159
        55600 => X"A8",  -- 168
        55601 => X"A4",  -- 164
        55602 => X"A5",  -- 165
        55603 => X"9E",  -- 158
        55604 => X"8E",  -- 142
        55605 => X"8A",  -- 138
        55606 => X"9A",  -- 154
        55607 => X"A5",  -- 165
        55608 => X"AA",  -- 170
        55609 => X"A0",  -- 160
        55610 => X"9D",  -- 157
        55611 => X"9F",  -- 159
        55612 => X"9F",  -- 159
        55613 => X"A3",  -- 163
        55614 => X"A6",  -- 166
        55615 => X"A5",  -- 165
        55616 => X"97",  -- 151
        55617 => X"8C",  -- 140
        55618 => X"8A",  -- 138
        55619 => X"99",  -- 153
        55620 => X"A6",  -- 166
        55621 => X"AC",  -- 172
        55622 => X"B1",  -- 177
        55623 => X"B8",  -- 184
        55624 => X"BD",  -- 189
        55625 => X"C3",  -- 195
        55626 => X"C8",  -- 200
        55627 => X"C8",  -- 200
        55628 => X"C5",  -- 197
        55629 => X"C5",  -- 197
        55630 => X"C7",  -- 199
        55631 => X"CC",  -- 204
        55632 => X"D0",  -- 208
        55633 => X"BC",  -- 188
        55634 => X"8B",  -- 139
        55635 => X"8D",  -- 141
        55636 => X"8E",  -- 142
        55637 => X"85",  -- 133
        55638 => X"80",  -- 128
        55639 => X"8D",  -- 141
        55640 => X"9F",  -- 159
        55641 => X"92",  -- 146
        55642 => X"8D",  -- 141
        55643 => X"8E",  -- 142
        55644 => X"8A",  -- 138
        55645 => X"8C",  -- 140
        55646 => X"8F",  -- 143
        55647 => X"89",  -- 137
        55648 => X"8D",  -- 141
        55649 => X"79",  -- 121
        55650 => X"61",  -- 97
        55651 => X"5E",  -- 94
        55652 => X"56",  -- 86
        55653 => X"4F",  -- 79
        55654 => X"4F",  -- 79
        55655 => X"3E",  -- 62
        55656 => X"49",  -- 73
        55657 => X"59",  -- 89
        55658 => X"45",  -- 69
        55659 => X"3E",  -- 62
        55660 => X"36",  -- 54
        55661 => X"36",  -- 54
        55662 => X"52",  -- 82
        55663 => X"4E",  -- 78
        55664 => X"42",  -- 66
        55665 => X"44",  -- 68
        55666 => X"4A",  -- 74
        55667 => X"4C",  -- 76
        55668 => X"4F",  -- 79
        55669 => X"56",  -- 86
        55670 => X"66",  -- 102
        55671 => X"75",  -- 117
        55672 => X"7C",  -- 124
        55673 => X"79",  -- 121
        55674 => X"67",  -- 103
        55675 => X"55",  -- 85
        55676 => X"50",  -- 80
        55677 => X"4E",  -- 78
        55678 => X"4A",  -- 74
        55679 => X"4D",  -- 77
        55680 => X"2D",  -- 45
        55681 => X"2D",  -- 45
        55682 => X"2C",  -- 44
        55683 => X"2C",  -- 44
        55684 => X"2B",  -- 43
        55685 => X"2C",  -- 44
        55686 => X"2C",  -- 44
        55687 => X"2C",  -- 44
        55688 => X"2E",  -- 46
        55689 => X"28",  -- 40
        55690 => X"25",  -- 37
        55691 => X"27",  -- 39
        55692 => X"2D",  -- 45
        55693 => X"2B",  -- 43
        55694 => X"23",  -- 35
        55695 => X"1B",  -- 27
        55696 => X"22",  -- 34
        55697 => X"38",  -- 56
        55698 => X"48",  -- 72
        55699 => X"3E",  -- 62
        55700 => X"2D",  -- 45
        55701 => X"23",  -- 35
        55702 => X"24",  -- 36
        55703 => X"27",  -- 39
        55704 => X"2B",  -- 43
        55705 => X"2F",  -- 47
        55706 => X"2F",  -- 47
        55707 => X"30",  -- 48
        55708 => X"35",  -- 53
        55709 => X"38",  -- 56
        55710 => X"31",  -- 49
        55711 => X"26",  -- 38
        55712 => X"22",  -- 34
        55713 => X"1D",  -- 29
        55714 => X"19",  -- 25
        55715 => X"19",  -- 25
        55716 => X"18",  -- 24
        55717 => X"1A",  -- 26
        55718 => X"22",  -- 34
        55719 => X"2A",  -- 42
        55720 => X"2B",  -- 43
        55721 => X"2C",  -- 44
        55722 => X"16",  -- 22
        55723 => X"25",  -- 37
        55724 => X"47",  -- 71
        55725 => X"24",  -- 36
        55726 => X"14",  -- 20
        55727 => X"4E",  -- 78
        55728 => X"4A",  -- 74
        55729 => X"3F",  -- 63
        55730 => X"2F",  -- 47
        55731 => X"21",  -- 33
        55732 => X"21",  -- 33
        55733 => X"2B",  -- 43
        55734 => X"31",  -- 49
        55735 => X"30",  -- 48
        55736 => X"26",  -- 38
        55737 => X"23",  -- 35
        55738 => X"5D",  -- 93
        55739 => X"8B",  -- 139
        55740 => X"63",  -- 99
        55741 => X"5C",  -- 92
        55742 => X"82",  -- 130
        55743 => X"72",  -- 114
        55744 => X"59",  -- 89
        55745 => X"54",  -- 84
        55746 => X"32",  -- 50
        55747 => X"18",  -- 24
        55748 => X"1F",  -- 31
        55749 => X"2A",  -- 42
        55750 => X"3C",  -- 60
        55751 => X"5B",  -- 91
        55752 => X"81",  -- 129
        55753 => X"A6",  -- 166
        55754 => X"A9",  -- 169
        55755 => X"91",  -- 145
        55756 => X"88",  -- 136
        55757 => X"77",  -- 119
        55758 => X"42",  -- 66
        55759 => X"10",  -- 16
        55760 => X"12",  -- 18
        55761 => X"1F",  -- 31
        55762 => X"32",  -- 50
        55763 => X"41",  -- 65
        55764 => X"46",  -- 70
        55765 => X"47",  -- 71
        55766 => X"4C",  -- 76
        55767 => X"53",  -- 83
        55768 => X"51",  -- 81
        55769 => X"59",  -- 89
        55770 => X"6A",  -- 106
        55771 => X"79",  -- 121
        55772 => X"74",  -- 116
        55773 => X"75",  -- 117
        55774 => X"70",  -- 112
        55775 => X"68",  -- 104
        55776 => X"66",  -- 102
        55777 => X"70",  -- 112
        55778 => X"6D",  -- 109
        55779 => X"5C",  -- 92
        55780 => X"4F",  -- 79
        55781 => X"4C",  -- 76
        55782 => X"48",  -- 72
        55783 => X"40",  -- 64
        55784 => X"38",  -- 56
        55785 => X"3B",  -- 59
        55786 => X"1D",  -- 29
        55787 => X"1C",  -- 28
        55788 => X"5A",  -- 90
        55789 => X"81",  -- 129
        55790 => X"BC",  -- 188
        55791 => X"D0",  -- 208
        55792 => X"D5",  -- 213
        55793 => X"BF",  -- 191
        55794 => X"90",  -- 144
        55795 => X"82",  -- 130
        55796 => X"73",  -- 115
        55797 => X"63",  -- 99
        55798 => X"5D",  -- 93
        55799 => X"2D",  -- 45
        55800 => X"56",  -- 86
        55801 => X"A5",  -- 165
        55802 => X"B5",  -- 181
        55803 => X"A5",  -- 165
        55804 => X"78",  -- 120
        55805 => X"85",  -- 133
        55806 => X"C8",  -- 200
        55807 => X"C8",  -- 200
        55808 => X"D2",  -- 210
        55809 => X"BA",  -- 186
        55810 => X"9B",  -- 155
        55811 => X"6E",  -- 110
        55812 => X"62",  -- 98
        55813 => X"53",  -- 83
        55814 => X"5A",  -- 90
        55815 => X"58",  -- 88
        55816 => X"4C",  -- 76
        55817 => X"51",  -- 81
        55818 => X"61",  -- 97
        55819 => X"71",  -- 113
        55820 => X"67",  -- 103
        55821 => X"64",  -- 100
        55822 => X"4F",  -- 79
        55823 => X"57",  -- 87
        55824 => X"44",  -- 68
        55825 => X"49",  -- 73
        55826 => X"52",  -- 82
        55827 => X"4A",  -- 74
        55828 => X"47",  -- 71
        55829 => X"5A",  -- 90
        55830 => X"49",  -- 73
        55831 => X"43",  -- 67
        55832 => X"33",  -- 51
        55833 => X"43",  -- 67
        55834 => X"53",  -- 83
        55835 => X"51",  -- 81
        55836 => X"45",  -- 69
        55837 => X"6F",  -- 111
        55838 => X"A0",  -- 160
        55839 => X"B1",  -- 177
        55840 => X"94",  -- 148
        55841 => X"87",  -- 135
        55842 => X"72",  -- 114
        55843 => X"52",  -- 82
        55844 => X"38",  -- 56
        55845 => X"41",  -- 65
        55846 => X"48",  -- 72
        55847 => X"3A",  -- 58
        55848 => X"1E",  -- 30
        55849 => X"1E",  -- 30
        55850 => X"1E",  -- 30
        55851 => X"25",  -- 37
        55852 => X"2D",  -- 45
        55853 => X"34",  -- 52
        55854 => X"38",  -- 56
        55855 => X"37",  -- 55
        55856 => X"34",  -- 52
        55857 => X"36",  -- 54
        55858 => X"36",  -- 54
        55859 => X"38",  -- 56
        55860 => X"3B",  -- 59
        55861 => X"3F",  -- 63
        55862 => X"46",  -- 70
        55863 => X"4A",  -- 74
        55864 => X"50",  -- 80
        55865 => X"4E",  -- 78
        55866 => X"4B",  -- 75
        55867 => X"4E",  -- 78
        55868 => X"57",  -- 87
        55869 => X"5F",  -- 95
        55870 => X"5D",  -- 93
        55871 => X"54",  -- 84
        55872 => X"4D",  -- 77
        55873 => X"50",  -- 80
        55874 => X"51",  -- 81
        55875 => X"51",  -- 81
        55876 => X"56",  -- 86
        55877 => X"61",  -- 97
        55878 => X"68",  -- 104
        55879 => X"6A",  -- 106
        55880 => X"68",  -- 104
        55881 => X"65",  -- 101
        55882 => X"60",  -- 96
        55883 => X"59",  -- 89
        55884 => X"4D",  -- 77
        55885 => X"44",  -- 68
        55886 => X"45",  -- 69
        55887 => X"4C",  -- 76
        55888 => X"47",  -- 71
        55889 => X"45",  -- 69
        55890 => X"45",  -- 69
        55891 => X"42",  -- 66
        55892 => X"40",  -- 64
        55893 => X"40",  -- 64
        55894 => X"41",  -- 65
        55895 => X"44",  -- 68
        55896 => X"6D",  -- 109
        55897 => X"80",  -- 128
        55898 => X"99",  -- 153
        55899 => X"AB",  -- 171
        55900 => X"B0",  -- 176
        55901 => X"AA",  -- 170
        55902 => X"A4",  -- 164
        55903 => X"A2",  -- 162
        55904 => X"A9",  -- 169
        55905 => X"A5",  -- 165
        55906 => X"A9",  -- 169
        55907 => X"AF",  -- 175
        55908 => X"AB",  -- 171
        55909 => X"9B",  -- 155
        55910 => X"92",  -- 146
        55911 => X"95",  -- 149
        55912 => X"93",  -- 147
        55913 => X"89",  -- 137
        55914 => X"93",  -- 147
        55915 => X"A2",  -- 162
        55916 => X"A4",  -- 164
        55917 => X"A6",  -- 166
        55918 => X"9D",  -- 157
        55919 => X"8F",  -- 143
        55920 => X"9D",  -- 157
        55921 => X"A8",  -- 168
        55922 => X"A9",  -- 169
        55923 => X"A2",  -- 162
        55924 => X"9E",  -- 158
        55925 => X"9C",  -- 156
        55926 => X"9F",  -- 159
        55927 => X"A5",  -- 165
        55928 => X"87",  -- 135
        55929 => X"8C",  -- 140
        55930 => X"8D",  -- 141
        55931 => X"8D",  -- 141
        55932 => X"86",  -- 134
        55933 => X"7D",  -- 125
        55934 => X"8A",  -- 138
        55935 => X"A6",  -- 166
        55936 => X"B1",  -- 177
        55937 => X"B2",  -- 178
        55938 => X"AA",  -- 170
        55939 => X"A0",  -- 160
        55940 => X"9E",  -- 158
        55941 => X"A8",  -- 168
        55942 => X"B4",  -- 180
        55943 => X"BA",  -- 186
        55944 => X"BC",  -- 188
        55945 => X"C1",  -- 193
        55946 => X"C4",  -- 196
        55947 => X"C5",  -- 197
        55948 => X"C5",  -- 197
        55949 => X"C6",  -- 198
        55950 => X"CC",  -- 204
        55951 => X"CF",  -- 207
        55952 => X"D3",  -- 211
        55953 => X"BC",  -- 188
        55954 => X"87",  -- 135
        55955 => X"8D",  -- 141
        55956 => X"8B",  -- 139
        55957 => X"80",  -- 128
        55958 => X"74",  -- 116
        55959 => X"82",  -- 130
        55960 => X"95",  -- 149
        55961 => X"91",  -- 145
        55962 => X"8E",  -- 142
        55963 => X"87",  -- 135
        55964 => X"7D",  -- 125
        55965 => X"81",  -- 129
        55966 => X"86",  -- 134
        55967 => X"7F",  -- 127
        55968 => X"83",  -- 131
        55969 => X"77",  -- 119
        55970 => X"62",  -- 98
        55971 => X"58",  -- 88
        55972 => X"48",  -- 72
        55973 => X"42",  -- 66
        55974 => X"4B",  -- 75
        55975 => X"42",  -- 66
        55976 => X"3D",  -- 61
        55977 => X"41",  -- 65
        55978 => X"3F",  -- 63
        55979 => X"3D",  -- 61
        55980 => X"3B",  -- 59
        55981 => X"3C",  -- 60
        55982 => X"46",  -- 70
        55983 => X"48",  -- 72
        55984 => X"51",  -- 81
        55985 => X"51",  -- 81
        55986 => X"53",  -- 83
        55987 => X"50",  -- 80
        55988 => X"4C",  -- 76
        55989 => X"4C",  -- 76
        55990 => X"5A",  -- 90
        55991 => X"69",  -- 105
        55992 => X"76",  -- 118
        55993 => X"73",  -- 115
        55994 => X"67",  -- 103
        55995 => X"5A",  -- 90
        55996 => X"50",  -- 80
        55997 => X"43",  -- 67
        55998 => X"42",  -- 66
        55999 => X"50",  -- 80
        56000 => X"25",  -- 37
        56001 => X"25",  -- 37
        56002 => X"26",  -- 38
        56003 => X"27",  -- 39
        56004 => X"27",  -- 39
        56005 => X"2B",  -- 43
        56006 => X"2C",  -- 44
        56007 => X"2E",  -- 46
        56008 => X"29",  -- 41
        56009 => X"23",  -- 35
        56010 => X"1F",  -- 31
        56011 => X"1F",  -- 31
        56012 => X"26",  -- 38
        56013 => X"2A",  -- 42
        56014 => X"29",  -- 41
        56015 => X"25",  -- 37
        56016 => X"2B",  -- 43
        56017 => X"3C",  -- 60
        56018 => X"43",  -- 67
        56019 => X"3A",  -- 58
        56020 => X"33",  -- 51
        56021 => X"33",  -- 51
        56022 => X"32",  -- 50
        56023 => X"29",  -- 41
        56024 => X"35",  -- 53
        56025 => X"2E",  -- 46
        56026 => X"2A",  -- 42
        56027 => X"2E",  -- 46
        56028 => X"32",  -- 50
        56029 => X"2D",  -- 45
        56030 => X"23",  -- 35
        56031 => X"1C",  -- 28
        56032 => X"19",  -- 25
        56033 => X"16",  -- 22
        56034 => X"14",  -- 20
        56035 => X"17",  -- 23
        56036 => X"1C",  -- 28
        56037 => X"20",  -- 32
        56038 => X"28",  -- 40
        56039 => X"33",  -- 51
        56040 => X"32",  -- 50
        56041 => X"1C",  -- 28
        56042 => X"2E",  -- 46
        56043 => X"3A",  -- 58
        56044 => X"1E",  -- 30
        56045 => X"27",  -- 39
        56046 => X"47",  -- 71
        56047 => X"47",  -- 71
        56048 => X"42",  -- 66
        56049 => X"2C",  -- 44
        56050 => X"22",  -- 34
        56051 => X"2F",  -- 47
        56052 => X"3A",  -- 58
        56053 => X"35",  -- 53
        56054 => X"31",  -- 49
        56055 => X"33",  -- 51
        56056 => X"42",  -- 66
        56057 => X"6A",  -- 106
        56058 => X"75",  -- 117
        56059 => X"6A",  -- 106
        56060 => X"63",  -- 99
        56061 => X"70",  -- 112
        56062 => X"78",  -- 120
        56063 => X"63",  -- 99
        56064 => X"6B",  -- 107
        56065 => X"6E",  -- 110
        56066 => X"50",  -- 80
        56067 => X"2E",  -- 46
        56068 => X"22",  -- 34
        56069 => X"1B",  -- 27
        56070 => X"28",  -- 40
        56071 => X"50",  -- 80
        56072 => X"7E",  -- 126
        56073 => X"89",  -- 137
        56074 => X"9B",  -- 155
        56075 => X"9C",  -- 156
        56076 => X"91",  -- 145
        56077 => X"83",  -- 131
        56078 => X"5F",  -- 95
        56079 => X"2D",  -- 45
        56080 => X"0D",  -- 13
        56081 => X"07",  -- 7
        56082 => X"0C",  -- 12
        56083 => X"22",  -- 34
        56084 => X"3A",  -- 58
        56085 => X"47",  -- 71
        56086 => X"4A",  -- 74
        56087 => X"4B",  -- 75
        56088 => X"4C",  -- 76
        56089 => X"31",  -- 49
        56090 => X"52",  -- 82
        56091 => X"62",  -- 98
        56092 => X"55",  -- 85
        56093 => X"46",  -- 70
        56094 => X"61",  -- 97
        56095 => X"5D",  -- 93
        56096 => X"4C",  -- 76
        56097 => X"5E",  -- 94
        56098 => X"62",  -- 98
        56099 => X"53",  -- 83
        56100 => X"48",  -- 72
        56101 => X"45",  -- 69
        56102 => X"39",  -- 57
        56103 => X"27",  -- 39
        56104 => X"11",  -- 17
        56105 => X"0B",  -- 11
        56106 => X"19",  -- 25
        56107 => X"5E",  -- 94
        56108 => X"A6",  -- 166
        56109 => X"AB",  -- 171
        56110 => X"CC",  -- 204
        56111 => X"CC",  -- 204
        56112 => X"C2",  -- 194
        56113 => X"B5",  -- 181
        56114 => X"91",  -- 145
        56115 => X"80",  -- 128
        56116 => X"50",  -- 80
        56117 => X"2F",  -- 47
        56118 => X"4E",  -- 78
        56119 => X"4D",  -- 77
        56120 => X"90",  -- 144
        56121 => X"B7",  -- 183
        56122 => X"CE",  -- 206
        56123 => X"AE",  -- 174
        56124 => X"4D",  -- 77
        56125 => X"6A",  -- 106
        56126 => X"BC",  -- 188
        56127 => X"C7",  -- 199
        56128 => X"B4",  -- 180
        56129 => X"AA",  -- 170
        56130 => X"9C",  -- 156
        56131 => X"6C",  -- 108
        56132 => X"49",  -- 73
        56133 => X"3F",  -- 63
        56134 => X"62",  -- 98
        56135 => X"79",  -- 121
        56136 => X"4C",  -- 76
        56137 => X"4A",  -- 74
        56138 => X"51",  -- 81
        56139 => X"5F",  -- 95
        56140 => X"57",  -- 87
        56141 => X"58",  -- 88
        56142 => X"41",  -- 65
        56143 => X"47",  -- 71
        56144 => X"34",  -- 52
        56145 => X"46",  -- 70
        56146 => X"40",  -- 64
        56147 => X"47",  -- 71
        56148 => X"3E",  -- 62
        56149 => X"53",  -- 83
        56150 => X"55",  -- 85
        56151 => X"43",  -- 67
        56152 => X"39",  -- 57
        56153 => X"53",  -- 83
        56154 => X"51",  -- 81
        56155 => X"5B",  -- 91
        56156 => X"52",  -- 82
        56157 => X"45",  -- 69
        56158 => X"3A",  -- 58
        56159 => X"61",  -- 97
        56160 => X"96",  -- 150
        56161 => X"5F",  -- 95
        56162 => X"5E",  -- 94
        56163 => X"93",  -- 147
        56164 => X"9A",  -- 154
        56165 => X"72",  -- 114
        56166 => X"4C",  -- 76
        56167 => X"39",  -- 57
        56168 => X"2A",  -- 42
        56169 => X"23",  -- 35
        56170 => X"1F",  -- 31
        56171 => X"25",  -- 37
        56172 => X"33",  -- 51
        56173 => X"3A",  -- 58
        56174 => X"3A",  -- 58
        56175 => X"34",  -- 52
        56176 => X"35",  -- 53
        56177 => X"36",  -- 54
        56178 => X"35",  -- 53
        56179 => X"34",  -- 52
        56180 => X"36",  -- 54
        56181 => X"3A",  -- 58
        56182 => X"41",  -- 65
        56183 => X"45",  -- 69
        56184 => X"51",  -- 81
        56185 => X"4E",  -- 78
        56186 => X"4B",  -- 75
        56187 => X"4E",  -- 78
        56188 => X"58",  -- 88
        56189 => X"61",  -- 97
        56190 => X"5D",  -- 93
        56191 => X"52",  -- 82
        56192 => X"4B",  -- 75
        56193 => X"4E",  -- 78
        56194 => X"52",  -- 82
        56195 => X"50",  -- 80
        56196 => X"52",  -- 82
        56197 => X"59",  -- 89
        56198 => X"5D",  -- 93
        56199 => X"5D",  -- 93
        56200 => X"59",  -- 89
        56201 => X"57",  -- 87
        56202 => X"54",  -- 84
        56203 => X"51",  -- 81
        56204 => X"4C",  -- 76
        56205 => X"44",  -- 68
        56206 => X"43",  -- 67
        56207 => X"47",  -- 71
        56208 => X"49",  -- 73
        56209 => X"4A",  -- 74
        56210 => X"4A",  -- 74
        56211 => X"4A",  -- 74
        56212 => X"4A",  -- 74
        56213 => X"49",  -- 73
        56214 => X"4B",  -- 75
        56215 => X"4E",  -- 78
        56216 => X"7D",  -- 125
        56217 => X"8C",  -- 140
        56218 => X"A8",  -- 168
        56219 => X"B4",  -- 180
        56220 => X"B4",  -- 180
        56221 => X"B2",  -- 178
        56222 => X"AD",  -- 173
        56223 => X"A1",  -- 161
        56224 => X"AF",  -- 175
        56225 => X"AB",  -- 171
        56226 => X"A7",  -- 167
        56227 => X"A5",  -- 165
        56228 => X"A2",  -- 162
        56229 => X"9F",  -- 159
        56230 => X"9B",  -- 155
        56231 => X"98",  -- 152
        56232 => X"9E",  -- 158
        56233 => X"98",  -- 152
        56234 => X"9D",  -- 157
        56235 => X"AB",  -- 171
        56236 => X"9C",  -- 156
        56237 => X"8B",  -- 139
        56238 => X"8E",  -- 142
        56239 => X"81",  -- 129
        56240 => X"97",  -- 151
        56241 => X"A2",  -- 162
        56242 => X"9C",  -- 156
        56243 => X"9A",  -- 154
        56244 => X"A9",  -- 169
        56245 => X"A7",  -- 167
        56246 => X"94",  -- 148
        56247 => X"89",  -- 137
        56248 => X"8C",  -- 140
        56249 => X"85",  -- 133
        56250 => X"7A",  -- 122
        56251 => X"7E",  -- 126
        56252 => X"83",  -- 131
        56253 => X"71",  -- 113
        56254 => X"6B",  -- 107
        56255 => X"7E",  -- 126
        56256 => X"98",  -- 152
        56257 => X"B3",  -- 179
        56258 => X"BD",  -- 189
        56259 => X"AE",  -- 174
        56260 => X"A5",  -- 165
        56261 => X"B0",  -- 176
        56262 => X"BA",  -- 186
        56263 => X"B6",  -- 182
        56264 => X"B8",  -- 184
        56265 => X"BA",  -- 186
        56266 => X"BD",  -- 189
        56267 => X"BF",  -- 191
        56268 => X"C2",  -- 194
        56269 => X"C8",  -- 200
        56270 => X"CF",  -- 207
        56271 => X"D4",  -- 212
        56272 => X"D6",  -- 214
        56273 => X"BC",  -- 188
        56274 => X"86",  -- 134
        56275 => X"8D",  -- 141
        56276 => X"88",  -- 136
        56277 => X"7B",  -- 123
        56278 => X"6B",  -- 107
        56279 => X"78",  -- 120
        56280 => X"85",  -- 133
        56281 => X"93",  -- 147
        56282 => X"99",  -- 153
        56283 => X"85",  -- 133
        56284 => X"6E",  -- 110
        56285 => X"72",  -- 114
        56286 => X"80",  -- 128
        56287 => X"7E",  -- 126
        56288 => X"70",  -- 112
        56289 => X"6D",  -- 109
        56290 => X"62",  -- 98
        56291 => X"58",  -- 88
        56292 => X"3F",  -- 63
        56293 => X"30",  -- 48
        56294 => X"3F",  -- 63
        56295 => X"40",  -- 64
        56296 => X"37",  -- 55
        56297 => X"36",  -- 54
        56298 => X"45",  -- 69
        56299 => X"36",  -- 54
        56300 => X"32",  -- 50
        56301 => X"3F",  -- 63
        56302 => X"3E",  -- 62
        56303 => X"4C",  -- 76
        56304 => X"57",  -- 87
        56305 => X"57",  -- 87
        56306 => X"57",  -- 87
        56307 => X"53",  -- 83
        56308 => X"4C",  -- 76
        56309 => X"4B",  -- 75
        56310 => X"57",  -- 87
        56311 => X"67",  -- 103
        56312 => X"72",  -- 114
        56313 => X"70",  -- 112
        56314 => X"6B",  -- 107
        56315 => X"66",  -- 102
        56316 => X"55",  -- 85
        56317 => X"3C",  -- 60
        56318 => X"3A",  -- 58
        56319 => X"53",  -- 83
        56320 => X"27",  -- 39
        56321 => X"28",  -- 40
        56322 => X"28",  -- 40
        56323 => X"27",  -- 39
        56324 => X"29",  -- 41
        56325 => X"2E",  -- 46
        56326 => X"2E",  -- 46
        56327 => X"2A",  -- 42
        56328 => X"26",  -- 38
        56329 => X"27",  -- 39
        56330 => X"22",  -- 34
        56331 => X"1D",  -- 29
        56332 => X"23",  -- 35
        56333 => X"2D",  -- 45
        56334 => X"2E",  -- 46
        56335 => X"26",  -- 38
        56336 => X"32",  -- 50
        56337 => X"3D",  -- 61
        56338 => X"3E",  -- 62
        56339 => X"34",  -- 52
        56340 => X"2F",  -- 47
        56341 => X"34",  -- 52
        56342 => X"35",  -- 53
        56343 => X"2F",  -- 47
        56344 => X"31",  -- 49
        56345 => X"2C",  -- 44
        56346 => X"27",  -- 39
        56347 => X"25",  -- 37
        56348 => X"25",  -- 37
        56349 => X"25",  -- 37
        56350 => X"22",  -- 34
        56351 => X"1F",  -- 31
        56352 => X"11",  -- 17
        56353 => X"1F",  -- 31
        56354 => X"14",  -- 20
        56355 => X"1D",  -- 29
        56356 => X"1E",  -- 30
        56357 => X"18",  -- 24
        56358 => X"28",  -- 40
        56359 => X"31",  -- 49
        56360 => X"2B",  -- 43
        56361 => X"2A",  -- 42
        56362 => X"2D",  -- 45
        56363 => X"20",  -- 32
        56364 => X"38",  -- 56
        56365 => X"5B",  -- 91
        56366 => X"2A",  -- 42
        56367 => X"41",  -- 65
        56368 => X"3F",  -- 63
        56369 => X"36",  -- 54
        56370 => X"33",  -- 51
        56371 => X"43",  -- 67
        56372 => X"3E",  -- 62
        56373 => X"40",  -- 64
        56374 => X"54",  -- 84
        56375 => X"69",  -- 105
        56376 => X"79",  -- 121
        56377 => X"79",  -- 121
        56378 => X"6D",  -- 109
        56379 => X"48",  -- 72
        56380 => X"79",  -- 121
        56381 => X"8B",  -- 139
        56382 => X"7E",  -- 126
        56383 => X"42",  -- 66
        56384 => X"49",  -- 73
        56385 => X"6C",  -- 108
        56386 => X"76",  -- 118
        56387 => X"5C",  -- 92
        56388 => X"41",  -- 65
        56389 => X"31",  -- 49
        56390 => X"28",  -- 40
        56391 => X"27",  -- 39
        56392 => X"43",  -- 67
        56393 => X"90",  -- 144
        56394 => X"AB",  -- 171
        56395 => X"9A",  -- 154
        56396 => X"9F",  -- 159
        56397 => X"91",  -- 145
        56398 => X"67",  -- 103
        56399 => X"56",  -- 86
        56400 => X"28",  -- 40
        56401 => X"18",  -- 24
        56402 => X"08",  -- 8
        56403 => X"07",  -- 7
        56404 => X"20",  -- 32
        56405 => X"3A",  -- 58
        56406 => X"43",  -- 67
        56407 => X"40",  -- 64
        56408 => X"40",  -- 64
        56409 => X"2E",  -- 46
        56410 => X"2D",  -- 45
        56411 => X"3B",  -- 59
        56412 => X"3A",  -- 58
        56413 => X"2F",  -- 47
        56414 => X"34",  -- 52
        56415 => X"49",  -- 73
        56416 => X"38",  -- 56
        56417 => X"3D",  -- 61
        56418 => X"49",  -- 73
        56419 => X"53",  -- 83
        56420 => X"49",  -- 73
        56421 => X"2D",  -- 45
        56422 => X"10",  -- 16
        56423 => X"02",  -- 2
        56424 => X"0F",  -- 15
        56425 => X"1A",  -- 26
        56426 => X"44",  -- 68
        56427 => X"90",  -- 144
        56428 => X"B0",  -- 176
        56429 => X"A1",  -- 161
        56430 => X"AA",  -- 170
        56431 => X"BD",  -- 189
        56432 => X"AB",  -- 171
        56433 => X"B1",  -- 177
        56434 => X"79",  -- 121
        56435 => X"6B",  -- 107
        56436 => X"4D",  -- 77
        56437 => X"41",  -- 65
        56438 => X"85",  -- 133
        56439 => X"88",  -- 136
        56440 => X"B0",  -- 176
        56441 => X"B5",  -- 181
        56442 => X"C9",  -- 201
        56443 => X"B9",  -- 185
        56444 => X"6D",  -- 109
        56445 => X"77",  -- 119
        56446 => X"BF",  -- 191
        56447 => X"AF",  -- 175
        56448 => X"B7",  -- 183
        56449 => X"D8",  -- 216
        56450 => X"BB",  -- 187
        56451 => X"67",  -- 103
        56452 => X"50",  -- 80
        56453 => X"48",  -- 72
        56454 => X"32",  -- 50
        56455 => X"55",  -- 85
        56456 => X"7D",  -- 125
        56457 => X"99",  -- 153
        56458 => X"80",  -- 128
        56459 => X"78",  -- 120
        56460 => X"4A",  -- 74
        56461 => X"3B",  -- 59
        56462 => X"52",  -- 82
        56463 => X"4C",  -- 76
        56464 => X"32",  -- 50
        56465 => X"20",  -- 32
        56466 => X"43",  -- 67
        56467 => X"45",  -- 69
        56468 => X"39",  -- 57
        56469 => X"57",  -- 87
        56470 => X"59",  -- 89
        56471 => X"42",  -- 66
        56472 => X"40",  -- 64
        56473 => X"49",  -- 73
        56474 => X"47",  -- 71
        56475 => X"58",  -- 88
        56476 => X"52",  -- 82
        56477 => X"3E",  -- 62
        56478 => X"47",  -- 71
        56479 => X"45",  -- 69
        56480 => X"4A",  -- 74
        56481 => X"73",  -- 115
        56482 => X"72",  -- 114
        56483 => X"4E",  -- 78
        56484 => X"47",  -- 71
        56485 => X"58",  -- 88
        56486 => X"6B",  -- 107
        56487 => X"7D",  -- 125
        56488 => X"63",  -- 99
        56489 => X"49",  -- 73
        56490 => X"31",  -- 49
        56491 => X"1F",  -- 31
        56492 => X"31",  -- 49
        56493 => X"46",  -- 70
        56494 => X"40",  -- 64
        56495 => X"3B",  -- 59
        56496 => X"38",  -- 56
        56497 => X"3B",  -- 59
        56498 => X"3B",  -- 59
        56499 => X"35",  -- 53
        56500 => X"33",  -- 51
        56501 => X"3A",  -- 58
        56502 => X"43",  -- 67
        56503 => X"47",  -- 71
        56504 => X"4E",  -- 78
        56505 => X"52",  -- 82
        56506 => X"53",  -- 83
        56507 => X"54",  -- 84
        56508 => X"5A",  -- 90
        56509 => X"5D",  -- 93
        56510 => X"57",  -- 87
        56511 => X"4F",  -- 79
        56512 => X"48",  -- 72
        56513 => X"4C",  -- 76
        56514 => X"4E",  -- 78
        56515 => X"4C",  -- 76
        56516 => X"50",  -- 80
        56517 => X"58",  -- 88
        56518 => X"60",  -- 96
        56519 => X"61",  -- 97
        56520 => X"62",  -- 98
        56521 => X"57",  -- 87
        56522 => X"4B",  -- 75
        56523 => X"41",  -- 65
        56524 => X"3F",  -- 63
        56525 => X"45",  -- 69
        56526 => X"4C",  -- 76
        56527 => X"53",  -- 83
        56528 => X"51",  -- 81
        56529 => X"50",  -- 80
        56530 => X"58",  -- 88
        56531 => X"51",  -- 81
        56532 => X"55",  -- 85
        56533 => X"50",  -- 80
        56534 => X"42",  -- 66
        56535 => X"5E",  -- 94
        56536 => X"82",  -- 130
        56537 => X"A1",  -- 161
        56538 => X"B5",  -- 181
        56539 => X"AD",  -- 173
        56540 => X"A5",  -- 165
        56541 => X"AC",  -- 172
        56542 => X"B5",  -- 181
        56543 => X"B8",  -- 184
        56544 => X"A9",  -- 169
        56545 => X"B3",  -- 179
        56546 => X"B4",  -- 180
        56547 => X"AD",  -- 173
        56548 => X"AA",  -- 170
        56549 => X"AF",  -- 175
        56550 => X"B1",  -- 177
        56551 => X"AE",  -- 174
        56552 => X"B8",  -- 184
        56553 => X"B5",  -- 181
        56554 => X"B4",  -- 180
        56555 => X"AA",  -- 170
        56556 => X"9B",  -- 155
        56557 => X"93",  -- 147
        56558 => X"8E",  -- 142
        56559 => X"82",  -- 130
        56560 => X"89",  -- 137
        56561 => X"97",  -- 151
        56562 => X"AF",  -- 175
        56563 => X"AE",  -- 174
        56564 => X"A0",  -- 160
        56565 => X"A4",  -- 164
        56566 => X"AB",  -- 171
        56567 => X"99",  -- 153
        56568 => X"9F",  -- 159
        56569 => X"9C",  -- 156
        56570 => X"98",  -- 152
        56571 => X"AA",  -- 170
        56572 => X"9F",  -- 159
        56573 => X"96",  -- 150
        56574 => X"77",  -- 119
        56575 => X"6D",  -- 109
        56576 => X"86",  -- 134
        56577 => X"A5",  -- 165
        56578 => X"C0",  -- 192
        56579 => X"C2",  -- 194
        56580 => X"B1",  -- 177
        56581 => X"B7",  -- 183
        56582 => X"C1",  -- 193
        56583 => X"AF",  -- 175
        56584 => X"B1",  -- 177
        56585 => X"B3",  -- 179
        56586 => X"B7",  -- 183
        56587 => X"B7",  -- 183
        56588 => X"BA",  -- 186
        56589 => X"C2",  -- 194
        56590 => X"CF",  -- 207
        56591 => X"DA",  -- 218
        56592 => X"DA",  -- 218
        56593 => X"B2",  -- 178
        56594 => X"7A",  -- 122
        56595 => X"75",  -- 117
        56596 => X"84",  -- 132
        56597 => X"7A",  -- 122
        56598 => X"6D",  -- 109
        56599 => X"6B",  -- 107
        56600 => X"73",  -- 115
        56601 => X"89",  -- 137
        56602 => X"8E",  -- 142
        56603 => X"88",  -- 136
        56604 => X"82",  -- 130
        56605 => X"6D",  -- 109
        56606 => X"60",  -- 96
        56607 => X"69",  -- 105
        56608 => X"67",  -- 103
        56609 => X"66",  -- 102
        56610 => X"5E",  -- 94
        56611 => X"52",  -- 82
        56612 => X"41",  -- 65
        56613 => X"2C",  -- 44
        56614 => X"27",  -- 39
        56615 => X"37",  -- 55
        56616 => X"39",  -- 57
        56617 => X"3B",  -- 59
        56618 => X"38",  -- 56
        56619 => X"32",  -- 50
        56620 => X"35",  -- 53
        56621 => X"40",  -- 64
        56622 => X"47",  -- 71
        56623 => X"46",  -- 70
        56624 => X"51",  -- 81
        56625 => X"53",  -- 83
        56626 => X"5C",  -- 92
        56627 => X"61",  -- 97
        56628 => X"55",  -- 85
        56629 => X"44",  -- 68
        56630 => X"4C",  -- 76
        56631 => X"62",  -- 98
        56632 => X"72",  -- 114
        56633 => X"73",  -- 115
        56634 => X"69",  -- 105
        56635 => X"5E",  -- 94
        56636 => X"59",  -- 89
        56637 => X"51",  -- 81
        56638 => X"4C",  -- 76
        56639 => X"53",  -- 83
        56640 => X"24",  -- 36
        56641 => X"25",  -- 37
        56642 => X"25",  -- 37
        56643 => X"24",  -- 36
        56644 => X"26",  -- 38
        56645 => X"2B",  -- 43
        56646 => X"2B",  -- 43
        56647 => X"27",  -- 39
        56648 => X"22",  -- 34
        56649 => X"23",  -- 35
        56650 => X"23",  -- 35
        56651 => X"1F",  -- 31
        56652 => X"1F",  -- 31
        56653 => X"24",  -- 36
        56654 => X"29",  -- 41
        56655 => X"2A",  -- 42
        56656 => X"32",  -- 50
        56657 => X"3B",  -- 59
        56658 => X"3B",  -- 59
        56659 => X"30",  -- 48
        56660 => X"2B",  -- 43
        56661 => X"30",  -- 48
        56662 => X"31",  -- 49
        56663 => X"2A",  -- 42
        56664 => X"2B",  -- 43
        56665 => X"27",  -- 39
        56666 => X"23",  -- 35
        56667 => X"21",  -- 33
        56668 => X"22",  -- 34
        56669 => X"23",  -- 35
        56670 => X"20",  -- 32
        56671 => X"1E",  -- 30
        56672 => X"1C",  -- 28
        56673 => X"11",  -- 17
        56674 => X"1E",  -- 30
        56675 => X"16",  -- 22
        56676 => X"25",  -- 37
        56677 => X"22",  -- 34
        56678 => X"1C",  -- 28
        56679 => X"28",  -- 40
        56680 => X"32",  -- 50
        56681 => X"20",  -- 32
        56682 => X"3E",  -- 62
        56683 => X"5C",  -- 92
        56684 => X"3B",  -- 59
        56685 => X"19",  -- 25
        56686 => X"4A",  -- 74
        56687 => X"5A",  -- 90
        56688 => X"5C",  -- 92
        56689 => X"3A",  -- 58
        56690 => X"39",  -- 57
        56691 => X"3D",  -- 61
        56692 => X"56",  -- 86
        56693 => X"6F",  -- 111
        56694 => X"64",  -- 100
        56695 => X"5E",  -- 94
        56696 => X"36",  -- 54
        56697 => X"52",  -- 82
        56698 => X"5D",  -- 93
        56699 => X"3E",  -- 62
        56700 => X"54",  -- 84
        56701 => X"5B",  -- 91
        56702 => X"57",  -- 87
        56703 => X"35",  -- 53
        56704 => X"38",  -- 56
        56705 => X"6D",  -- 109
        56706 => X"8B",  -- 139
        56707 => X"7F",  -- 127
        56708 => X"69",  -- 105
        56709 => X"52",  -- 82
        56710 => X"38",  -- 56
        56711 => X"26",  -- 38
        56712 => X"30",  -- 48
        56713 => X"69",  -- 105
        56714 => X"99",  -- 153
        56715 => X"A3",  -- 163
        56716 => X"9E",  -- 158
        56717 => X"94",  -- 148
        56718 => X"75",  -- 117
        56719 => X"4F",  -- 79
        56720 => X"48",  -- 72
        56721 => X"31",  -- 49
        56722 => X"18",  -- 24
        56723 => X"10",  -- 16
        56724 => X"14",  -- 20
        56725 => X"1D",  -- 29
        56726 => X"2D",  -- 45
        56727 => X"3A",  -- 58
        56728 => X"3C",  -- 60
        56729 => X"3A",  -- 58
        56730 => X"37",  -- 55
        56731 => X"31",  -- 49
        56732 => X"2C",  -- 44
        56733 => X"2B",  -- 43
        56734 => X"2D",  -- 45
        56735 => X"2D",  -- 45
        56736 => X"2D",  -- 45
        56737 => X"37",  -- 55
        56738 => X"43",  -- 67
        56739 => X"3D",  -- 61
        56740 => X"22",  -- 34
        56741 => X"0C",  -- 12
        56742 => X"10",  -- 16
        56743 => X"22",  -- 34
        56744 => X"3E",  -- 62
        56745 => X"64",  -- 100
        56746 => X"79",  -- 121
        56747 => X"89",  -- 137
        56748 => X"9E",  -- 158
        56749 => X"B9",  -- 185
        56750 => X"C5",  -- 197
        56751 => X"B1",  -- 177
        56752 => X"97",  -- 151
        56753 => X"5D",  -- 93
        56754 => X"35",  -- 53
        56755 => X"56",  -- 86
        56756 => X"71",  -- 113
        56757 => X"7A",  -- 122
        56758 => X"9E",  -- 158
        56759 => X"B3",  -- 179
        56760 => X"AA",  -- 170
        56761 => X"C5",  -- 197
        56762 => X"C3",  -- 195
        56763 => X"B4",  -- 180
        56764 => X"B4",  -- 180
        56765 => X"BD",  -- 189
        56766 => X"A9",  -- 169
        56767 => X"72",  -- 114
        56768 => X"A2",  -- 162
        56769 => X"CC",  -- 204
        56770 => X"B2",  -- 178
        56771 => X"64",  -- 100
        56772 => X"32",  -- 50
        56773 => X"2E",  -- 46
        56774 => X"40",  -- 64
        56775 => X"48",  -- 72
        56776 => X"40",  -- 64
        56777 => X"50",  -- 80
        56778 => X"84",  -- 132
        56779 => X"9F",  -- 159
        56780 => X"75",  -- 117
        56781 => X"55",  -- 85
        56782 => X"37",  -- 55
        56783 => X"4F",  -- 79
        56784 => X"95",  -- 149
        56785 => X"8E",  -- 142
        56786 => X"5A",  -- 90
        56787 => X"42",  -- 66
        56788 => X"2A",  -- 42
        56789 => X"51",  -- 81
        56790 => X"44",  -- 68
        56791 => X"55",  -- 85
        56792 => X"49",  -- 73
        56793 => X"47",  -- 71
        56794 => X"41",  -- 65
        56795 => X"53",  -- 83
        56796 => X"58",  -- 88
        56797 => X"49",  -- 73
        56798 => X"4A",  -- 74
        56799 => X"45",  -- 69
        56800 => X"48",  -- 72
        56801 => X"2B",  -- 43
        56802 => X"59",  -- 89
        56803 => X"86",  -- 134
        56804 => X"57",  -- 87
        56805 => X"2E",  -- 46
        56806 => X"35",  -- 53
        56807 => X"36",  -- 54
        56808 => X"24",  -- 36
        56809 => X"5D",  -- 93
        56810 => X"86",  -- 134
        56811 => X"6A",  -- 106
        56812 => X"51",  -- 81
        56813 => X"51",  -- 81
        56814 => X"45",  -- 69
        56815 => X"38",  -- 56
        56816 => X"45",  -- 69
        56817 => X"3C",  -- 60
        56818 => X"32",  -- 50
        56819 => X"2D",  -- 45
        56820 => X"2D",  -- 45
        56821 => X"34",  -- 52
        56822 => X"3F",  -- 63
        56823 => X"45",  -- 69
        56824 => X"48",  -- 72
        56825 => X"4E",  -- 78
        56826 => X"51",  -- 81
        56827 => X"51",  -- 81
        56828 => X"52",  -- 82
        56829 => X"52",  -- 82
        56830 => X"50",  -- 80
        56831 => X"4A",  -- 74
        56832 => X"5A",  -- 90
        56833 => X"57",  -- 87
        56834 => X"4D",  -- 77
        56835 => X"44",  -- 68
        56836 => X"43",  -- 67
        56837 => X"50",  -- 80
        56838 => X"61",  -- 97
        56839 => X"6B",  -- 107
        56840 => X"66",  -- 102
        56841 => X"5F",  -- 95
        56842 => X"56",  -- 86
        56843 => X"50",  -- 80
        56844 => X"51",  -- 81
        56845 => X"55",  -- 85
        56846 => X"5D",  -- 93
        56847 => X"60",  -- 96
        56848 => X"63",  -- 99
        56849 => X"5F",  -- 95
        56850 => X"61",  -- 97
        56851 => X"58",  -- 88
        56852 => X"57",  -- 87
        56853 => X"50",  -- 80
        56854 => X"4A",  -- 74
        56855 => X"6A",  -- 106
        56856 => X"90",  -- 144
        56857 => X"9A",  -- 154
        56858 => X"A2",  -- 162
        56859 => X"A4",  -- 164
        56860 => X"A9",  -- 169
        56861 => X"AE",  -- 174
        56862 => X"A6",  -- 166
        56863 => X"95",  -- 149
        56864 => X"A2",  -- 162
        56865 => X"B0",  -- 176
        56866 => X"BA",  -- 186
        56867 => X"B6",  -- 182
        56868 => X"B2",  -- 178
        56869 => X"B5",  -- 181
        56870 => X"B4",  -- 180
        56871 => X"B2",  -- 178
        56872 => X"B1",  -- 177
        56873 => X"AF",  -- 175
        56874 => X"B3",  -- 179
        56875 => X"B2",  -- 178
        56876 => X"AA",  -- 170
        56877 => X"A7",  -- 167
        56878 => X"A1",  -- 161
        56879 => X"93",  -- 147
        56880 => X"7C",  -- 124
        56881 => X"9F",  -- 159
        56882 => X"C2",  -- 194
        56883 => X"C6",  -- 198
        56884 => X"A8",  -- 168
        56885 => X"AA",  -- 170
        56886 => X"B5",  -- 181
        56887 => X"B6",  -- 182
        56888 => X"C3",  -- 195
        56889 => X"BF",  -- 191
        56890 => X"B7",  -- 183
        56891 => X"BC",  -- 188
        56892 => X"B5",  -- 181
        56893 => X"AD",  -- 173
        56894 => X"99",  -- 153
        56895 => X"8F",  -- 143
        56896 => X"7D",  -- 125
        56897 => X"9A",  -- 154
        56898 => X"BA",  -- 186
        56899 => X"C2",  -- 194
        56900 => X"B7",  -- 183
        56901 => X"B4",  -- 180
        56902 => X"BD",  -- 189
        56903 => X"BD",  -- 189
        56904 => X"B7",  -- 183
        56905 => X"B6",  -- 182
        56906 => X"B5",  -- 181
        56907 => X"B3",  -- 179
        56908 => X"B3",  -- 179
        56909 => X"B9",  -- 185
        56910 => X"C1",  -- 193
        56911 => X"C9",  -- 201
        56912 => X"D7",  -- 215
        56913 => X"AF",  -- 175
        56914 => X"75",  -- 117
        56915 => X"72",  -- 114
        56916 => X"7F",  -- 127
        56917 => X"78",  -- 120
        56918 => X"6D",  -- 109
        56919 => X"4F",  -- 79
        56920 => X"61",  -- 97
        56921 => X"78",  -- 120
        56922 => X"86",  -- 134
        56923 => X"84",  -- 132
        56924 => X"7A",  -- 122
        56925 => X"68",  -- 104
        56926 => X"56",  -- 86
        56927 => X"4C",  -- 76
        56928 => X"55",  -- 85
        56929 => X"56",  -- 86
        56930 => X"51",  -- 81
        56931 => X"4B",  -- 75
        56932 => X"42",  -- 66
        56933 => X"30",  -- 48
        56934 => X"28",  -- 40
        56935 => X"32",  -- 50
        56936 => X"32",  -- 50
        56937 => X"35",  -- 53
        56938 => X"37",  -- 55
        56939 => X"36",  -- 54
        56940 => X"39",  -- 57
        56941 => X"3F",  -- 63
        56942 => X"43",  -- 67
        56943 => X"43",  -- 67
        56944 => X"4C",  -- 76
        56945 => X"4F",  -- 79
        56946 => X"5A",  -- 90
        56947 => X"63",  -- 99
        56948 => X"5F",  -- 95
        56949 => X"50",  -- 80
        56950 => X"44",  -- 68
        56951 => X"42",  -- 66
        56952 => X"5E",  -- 94
        56953 => X"6D",  -- 109
        56954 => X"6D",  -- 109
        56955 => X"62",  -- 98
        56956 => X"5F",  -- 95
        56957 => X"5C",  -- 92
        56958 => X"5C",  -- 92
        56959 => X"5F",  -- 95
        56960 => X"23",  -- 35
        56961 => X"25",  -- 37
        56962 => X"24",  -- 36
        56963 => X"22",  -- 34
        56964 => X"24",  -- 36
        56965 => X"28",  -- 40
        56966 => X"27",  -- 39
        56967 => X"24",  -- 36
        56968 => X"1E",  -- 30
        56969 => X"20",  -- 32
        56970 => X"22",  -- 34
        56971 => X"20",  -- 32
        56972 => X"1E",  -- 30
        56973 => X"1E",  -- 30
        56974 => X"26",  -- 38
        56975 => X"31",  -- 49
        56976 => X"39",  -- 57
        56977 => X"3F",  -- 63
        56978 => X"3D",  -- 61
        56979 => X"31",  -- 49
        56980 => X"2C",  -- 44
        56981 => X"30",  -- 48
        56982 => X"2E",  -- 46
        56983 => X"25",  -- 37
        56984 => X"21",  -- 33
        56985 => X"1F",  -- 31
        56986 => X"1C",  -- 28
        56987 => X"1E",  -- 30
        56988 => X"21",  -- 33
        56989 => X"22",  -- 34
        56990 => X"21",  -- 33
        56991 => X"1F",  -- 31
        56992 => X"19",  -- 25
        56993 => X"1E",  -- 30
        56994 => X"1C",  -- 28
        56995 => X"1D",  -- 29
        56996 => X"22",  -- 34
        56997 => X"2A",  -- 42
        56998 => X"31",  -- 49
        56999 => X"30",  -- 48
        57000 => X"2D",  -- 45
        57001 => X"44",  -- 68
        57002 => X"64",  -- 100
        57003 => X"36",  -- 54
        57004 => X"2F",  -- 47
        57005 => X"77",  -- 119
        57006 => X"7D",  -- 125
        57007 => X"70",  -- 112
        57008 => X"52",  -- 82
        57009 => X"41",  -- 65
        57010 => X"4B",  -- 75
        57011 => X"77",  -- 119
        57012 => X"6C",  -- 108
        57013 => X"4E",  -- 78
        57014 => X"53",  -- 83
        57015 => X"2A",  -- 42
        57016 => X"27",  -- 39
        57017 => X"46",  -- 70
        57018 => X"5A",  -- 90
        57019 => X"4A",  -- 74
        57020 => X"40",  -- 64
        57021 => X"38",  -- 56
        57022 => X"4B",  -- 75
        57023 => X"60",  -- 96
        57024 => X"4F",  -- 79
        57025 => X"75",  -- 117
        57026 => X"88",  -- 136
        57027 => X"82",  -- 130
        57028 => X"81",  -- 129
        57029 => X"7B",  -- 123
        57030 => X"62",  -- 98
        57031 => X"48",  -- 72
        57032 => X"35",  -- 53
        57033 => X"4F",  -- 79
        57034 => X"87",  -- 135
        57035 => X"A0",  -- 160
        57036 => X"93",  -- 147
        57037 => X"99",  -- 153
        57038 => X"99",  -- 153
        57039 => X"77",  -- 119
        57040 => X"6E",  -- 110
        57041 => X"53",  -- 83
        57042 => X"3A",  -- 58
        57043 => X"2E",  -- 46
        57044 => X"1B",  -- 27
        57045 => X"0C",  -- 12
        57046 => X"14",  -- 20
        57047 => X"2B",  -- 43
        57048 => X"2C",  -- 44
        57049 => X"33",  -- 51
        57050 => X"32",  -- 50
        57051 => X"29",  -- 41
        57052 => X"28",  -- 40
        57053 => X"2E",  -- 46
        57054 => X"2C",  -- 44
        57055 => X"25",  -- 37
        57056 => X"31",  -- 49
        57057 => X"38",  -- 56
        57058 => X"31",  -- 49
        57059 => X"1D",  -- 29
        57060 => X"0F",  -- 15
        57061 => X"1C",  -- 28
        57062 => X"36",  -- 54
        57063 => X"49",  -- 73
        57064 => X"57",  -- 87
        57065 => X"7D",  -- 125
        57066 => X"94",  -- 148
        57067 => X"AA",  -- 170
        57068 => X"BF",  -- 191
        57069 => X"CC",  -- 204
        57070 => X"CB",  -- 203
        57071 => X"AF",  -- 175
        57072 => X"85",  -- 133
        57073 => X"45",  -- 69
        57074 => X"4D",  -- 77
        57075 => X"7B",  -- 123
        57076 => X"9D",  -- 157
        57077 => X"A6",  -- 166
        57078 => X"A7",  -- 167
        57079 => X"CB",  -- 203
        57080 => X"BF",  -- 191
        57081 => X"A6",  -- 166
        57082 => X"BA",  -- 186
        57083 => X"CC",  -- 204
        57084 => X"B5",  -- 181
        57085 => X"9C",  -- 156
        57086 => X"96",  -- 150
        57087 => X"A2",  -- 162
        57088 => X"B8",  -- 184
        57089 => X"A7",  -- 167
        57090 => X"97",  -- 151
        57091 => X"8B",  -- 139
        57092 => X"4F",  -- 79
        57093 => X"39",  -- 57
        57094 => X"56",  -- 86
        57095 => X"37",  -- 55
        57096 => X"3D",  -- 61
        57097 => X"3B",  -- 59
        57098 => X"27",  -- 39
        57099 => X"5C",  -- 92
        57100 => X"61",  -- 97
        57101 => X"6E",  -- 110
        57102 => X"73",  -- 115
        57103 => X"25",  -- 37
        57104 => X"3C",  -- 60
        57105 => X"55",  -- 85
        57106 => X"93",  -- 147
        57107 => X"A2",  -- 162
        57108 => X"7E",  -- 126
        57109 => X"5E",  -- 94
        57110 => X"67",  -- 103
        57111 => X"4A",  -- 74
        57112 => X"3E",  -- 62
        57113 => X"4B",  -- 75
        57114 => X"49",  -- 73
        57115 => X"45",  -- 69
        57116 => X"43",  -- 67
        57117 => X"46",  -- 70
        57118 => X"50",  -- 80
        57119 => X"4B",  -- 75
        57120 => X"3E",  -- 62
        57121 => X"47",  -- 71
        57122 => X"29",  -- 41
        57123 => X"36",  -- 54
        57124 => X"72",  -- 114
        57125 => X"62",  -- 98
        57126 => X"20",  -- 32
        57127 => X"15",  -- 21
        57128 => X"33",  -- 51
        57129 => X"09",  -- 9
        57130 => X"17",  -- 23
        57131 => X"43",  -- 67
        57132 => X"68",  -- 104
        57133 => X"88",  -- 136
        57134 => X"7B",  -- 123
        57135 => X"5B",  -- 91
        57136 => X"49",  -- 73
        57137 => X"3F",  -- 63
        57138 => X"39",  -- 57
        57139 => X"3B",  -- 59
        57140 => X"3E",  -- 62
        57141 => X"3D",  -- 61
        57142 => X"3F",  -- 63
        57143 => X"45",  -- 69
        57144 => X"44",  -- 68
        57145 => X"48",  -- 72
        57146 => X"4A",  -- 74
        57147 => X"46",  -- 70
        57148 => X"42",  -- 66
        57149 => X"42",  -- 66
        57150 => X"41",  -- 65
        57151 => X"42",  -- 66
        57152 => X"42",  -- 66
        57153 => X"4A",  -- 74
        57154 => X"4F",  -- 79
        57155 => X"52",  -- 82
        57156 => X"54",  -- 84
        57157 => X"5C",  -- 92
        57158 => X"66",  -- 102
        57159 => X"6C",  -- 108
        57160 => X"6E",  -- 110
        57161 => X"6B",  -- 107
        57162 => X"66",  -- 102
        57163 => X"65",  -- 101
        57164 => X"65",  -- 101
        57165 => X"69",  -- 105
        57166 => X"6D",  -- 109
        57167 => X"6F",  -- 111
        57168 => X"6E",  -- 110
        57169 => X"63",  -- 99
        57170 => X"60",  -- 96
        57171 => X"57",  -- 87
        57172 => X"50",  -- 80
        57173 => X"4B",  -- 75
        57174 => X"55",  -- 85
        57175 => X"7C",  -- 124
        57176 => X"96",  -- 150
        57177 => X"95",  -- 149
        57178 => X"94",  -- 148
        57179 => X"92",  -- 146
        57180 => X"95",  -- 149
        57181 => X"97",  -- 151
        57182 => X"95",  -- 149
        57183 => X"90",  -- 144
        57184 => X"A1",  -- 161
        57185 => X"AE",  -- 174
        57186 => X"B9",  -- 185
        57187 => X"BA",  -- 186
        57188 => X"B7",  -- 183
        57189 => X"B7",  -- 183
        57190 => X"B9",  -- 185
        57191 => X"B7",  -- 183
        57192 => X"AB",  -- 171
        57193 => X"A9",  -- 169
        57194 => X"AC",  -- 172
        57195 => X"AD",  -- 173
        57196 => X"A7",  -- 167
        57197 => X"A8",  -- 168
        57198 => X"A4",  -- 164
        57199 => X"98",  -- 152
        57200 => X"9A",  -- 154
        57201 => X"B2",  -- 178
        57202 => X"BC",  -- 188
        57203 => X"BD",  -- 189
        57204 => X"98",  -- 152
        57205 => X"A5",  -- 165
        57206 => X"AA",  -- 170
        57207 => X"B2",  -- 178
        57208 => X"AC",  -- 172
        57209 => X"B0",  -- 176
        57210 => X"BB",  -- 187
        57211 => X"BC",  -- 188
        57212 => X"C6",  -- 198
        57213 => X"C5",  -- 197
        57214 => X"C2",  -- 194
        57215 => X"B8",  -- 184
        57216 => X"97",  -- 151
        57217 => X"A7",  -- 167
        57218 => X"B7",  -- 183
        57219 => X"BC",  -- 188
        57220 => X"B8",  -- 184
        57221 => X"AD",  -- 173
        57222 => X"AA",  -- 170
        57223 => X"B6",  -- 182
        57224 => X"B3",  -- 179
        57225 => X"B3",  -- 179
        57226 => X"B4",  -- 180
        57227 => X"B5",  -- 181
        57228 => X"B7",  -- 183
        57229 => X"B9",  -- 185
        57230 => X"BB",  -- 187
        57231 => X"BD",  -- 189
        57232 => X"D6",  -- 214
        57233 => X"B4",  -- 180
        57234 => X"6F",  -- 111
        57235 => X"65",  -- 101
        57236 => X"6E",  -- 110
        57237 => X"70",  -- 112
        57238 => X"7D",  -- 125
        57239 => X"5D",  -- 93
        57240 => X"4C",  -- 76
        57241 => X"5B",  -- 91
        57242 => X"70",  -- 112
        57243 => X"79",  -- 121
        57244 => X"70",  -- 112
        57245 => X"64",  -- 100
        57246 => X"53",  -- 83
        57247 => X"3E",  -- 62
        57248 => X"3F",  -- 63
        57249 => X"40",  -- 64
        57250 => X"3D",  -- 61
        57251 => X"3F",  -- 63
        57252 => X"41",  -- 65
        57253 => X"34",  -- 52
        57254 => X"29",  -- 41
        57255 => X"2D",  -- 45
        57256 => X"2F",  -- 47
        57257 => X"2F",  -- 47
        57258 => X"32",  -- 50
        57259 => X"37",  -- 55
        57260 => X"39",  -- 57
        57261 => X"3B",  -- 59
        57262 => X"41",  -- 65
        57263 => X"47",  -- 71
        57264 => X"42",  -- 66
        57265 => X"49",  -- 73
        57266 => X"52",  -- 82
        57267 => X"5C",  -- 92
        57268 => X"66",  -- 102
        57269 => X"64",  -- 100
        57270 => X"50",  -- 80
        57271 => X"39",  -- 57
        57272 => X"43",  -- 67
        57273 => X"5D",  -- 93
        57274 => X"66",  -- 102
        57275 => X"5E",  -- 94
        57276 => X"5D",  -- 93
        57277 => X"60",  -- 96
        57278 => X"64",  -- 100
        57279 => X"69",  -- 105
        57280 => X"26",  -- 38
        57281 => X"27",  -- 39
        57282 => X"25",  -- 37
        57283 => X"23",  -- 35
        57284 => X"24",  -- 36
        57285 => X"27",  -- 39
        57286 => X"25",  -- 37
        57287 => X"21",  -- 33
        57288 => X"1E",  -- 30
        57289 => X"1C",  -- 28
        57290 => X"1E",  -- 30
        57291 => X"22",  -- 34
        57292 => X"20",  -- 32
        57293 => X"1D",  -- 29
        57294 => X"26",  -- 38
        57295 => X"33",  -- 51
        57296 => X"43",  -- 67
        57297 => X"47",  -- 71
        57298 => X"43",  -- 67
        57299 => X"36",  -- 54
        57300 => X"31",  -- 49
        57301 => X"31",  -- 49
        57302 => X"2C",  -- 44
        57303 => X"24",  -- 36
        57304 => X"1C",  -- 28
        57305 => X"1A",  -- 26
        57306 => X"1B",  -- 27
        57307 => X"1C",  -- 28
        57308 => X"20",  -- 32
        57309 => X"24",  -- 36
        57310 => X"25",  -- 37
        57311 => X"25",  -- 37
        57312 => X"24",  -- 36
        57313 => X"25",  -- 37
        57314 => X"17",  -- 23
        57315 => X"1A",  -- 26
        57316 => X"0D",  -- 13
        57317 => X"31",  -- 49
        57318 => X"20",  -- 32
        57319 => X"18",  -- 24
        57320 => X"54",  -- 84
        57321 => X"8E",  -- 142
        57322 => X"5C",  -- 92
        57323 => X"6A",  -- 106
        57324 => X"68",  -- 104
        57325 => X"7D",  -- 125
        57326 => X"55",  -- 85
        57327 => X"47",  -- 71
        57328 => X"39",  -- 57
        57329 => X"6B",  -- 107
        57330 => X"7F",  -- 127
        57331 => X"34",  -- 52
        57332 => X"2C",  -- 44
        57333 => X"3E",  -- 62
        57334 => X"33",  -- 51
        57335 => X"46",  -- 70
        57336 => X"66",  -- 102
        57337 => X"58",  -- 88
        57338 => X"51",  -- 81
        57339 => X"61",  -- 97
        57340 => X"60",  -- 96
        57341 => X"43",  -- 67
        57342 => X"2F",  -- 47
        57343 => X"39",  -- 57
        57344 => X"5C",  -- 92
        57345 => X"74",  -- 116
        57346 => X"81",  -- 129
        57347 => X"82",  -- 130
        57348 => X"86",  -- 134
        57349 => X"82",  -- 130
        57350 => X"72",  -- 114
        57351 => X"68",  -- 104
        57352 => X"5F",  -- 95
        57353 => X"61",  -- 97
        57354 => X"7F",  -- 127
        57355 => X"90",  -- 144
        57356 => X"85",  -- 133
        57357 => X"90",  -- 144
        57358 => X"9D",  -- 157
        57359 => X"8D",  -- 141
        57360 => X"82",  -- 130
        57361 => X"71",  -- 113
        57362 => X"62",  -- 98
        57363 => X"55",  -- 85
        57364 => X"3B",  -- 59
        57365 => X"19",  -- 25
        57366 => X"0C",  -- 12
        57367 => X"13",  -- 19
        57368 => X"1C",  -- 28
        57369 => X"1B",  -- 27
        57370 => X"21",  -- 33
        57371 => X"27",  -- 39
        57372 => X"29",  -- 41
        57373 => X"28",  -- 40
        57374 => X"28",  -- 40
        57375 => X"2A",  -- 42
        57376 => X"2D",  -- 45
        57377 => X"30",  -- 48
        57378 => X"1D",  -- 29
        57379 => X"09",  -- 9
        57380 => X"1A",  -- 26
        57381 => X"4D",  -- 77
        57382 => X"6B",  -- 107
        57383 => X"6B",  -- 107
        57384 => X"81",  -- 129
        57385 => X"8B",  -- 139
        57386 => X"97",  -- 151
        57387 => X"B9",  -- 185
        57388 => X"CA",  -- 202
        57389 => X"C3",  -- 195
        57390 => X"C5",  -- 197
        57391 => X"C2",  -- 194
        57392 => X"A3",  -- 163
        57393 => X"81",  -- 129
        57394 => X"8F",  -- 143
        57395 => X"A3",  -- 163
        57396 => X"B9",  -- 185
        57397 => X"C4",  -- 196
        57398 => X"B0",  -- 176
        57399 => X"B0",  -- 176
        57400 => X"D3",  -- 211
        57401 => X"BB",  -- 187
        57402 => X"B5",  -- 181
        57403 => X"8C",  -- 140
        57404 => X"6C",  -- 108
        57405 => X"75",  -- 117
        57406 => X"73",  -- 115
        57407 => X"73",  -- 115
        57408 => X"B4",  -- 180
        57409 => X"97",  -- 151
        57410 => X"5E",  -- 94
        57411 => X"78",  -- 120
        57412 => X"AF",  -- 175
        57413 => X"8F",  -- 143
        57414 => X"59",  -- 89
        57415 => X"48",  -- 72
        57416 => X"2C",  -- 44
        57417 => X"43",  -- 67
        57418 => X"2D",  -- 45
        57419 => X"23",  -- 35
        57420 => X"32",  -- 50
        57421 => X"40",  -- 64
        57422 => X"41",  -- 65
        57423 => X"80",  -- 128
        57424 => X"56",  -- 86
        57425 => X"2E",  -- 46
        57426 => X"27",  -- 39
        57427 => X"39",  -- 57
        57428 => X"84",  -- 132
        57429 => X"88",  -- 136
        57430 => X"A2",  -- 162
        57431 => X"79",  -- 121
        57432 => X"5A",  -- 90
        57433 => X"43",  -- 67
        57434 => X"3B",  -- 59
        57435 => X"51",  -- 81
        57436 => X"56",  -- 86
        57437 => X"44",  -- 68
        57438 => X"40",  -- 64
        57439 => X"4B",  -- 75
        57440 => X"4D",  -- 77
        57441 => X"3D",  -- 61
        57442 => X"3C",  -- 60
        57443 => X"2C",  -- 44
        57444 => X"22",  -- 34
        57445 => X"53",  -- 83
        57446 => X"66",  -- 102
        57447 => X"32",  -- 50
        57448 => X"06",  -- 6
        57449 => X"26",  -- 38
        57450 => X"2C",  -- 44
        57451 => X"21",  -- 33
        57452 => X"3C",  -- 60
        57453 => X"43",  -- 67
        57454 => X"3E",  -- 62
        57455 => X"5F",  -- 95
        57456 => X"82",  -- 130
        57457 => X"6D",  -- 109
        57458 => X"57",  -- 87
        57459 => X"4D",  -- 77
        57460 => X"45",  -- 69
        57461 => X"3C",  -- 60
        57462 => X"3D",  -- 61
        57463 => X"46",  -- 70
        57464 => X"45",  -- 69
        57465 => X"45",  -- 69
        57466 => X"40",  -- 64
        57467 => X"39",  -- 57
        57468 => X"32",  -- 50
        57469 => X"30",  -- 48
        57470 => X"33",  -- 51
        57471 => X"34",  -- 52
        57472 => X"40",  -- 64
        57473 => X"43",  -- 67
        57474 => X"44",  -- 68
        57475 => X"42",  -- 66
        57476 => X"47",  -- 71
        57477 => X"53",  -- 83
        57478 => X"65",  -- 101
        57479 => X"70",  -- 112
        57480 => X"77",  -- 119
        57481 => X"74",  -- 116
        57482 => X"73",  -- 115
        57483 => X"71",  -- 113
        57484 => X"71",  -- 113
        57485 => X"72",  -- 114
        57486 => X"71",  -- 113
        57487 => X"6F",  -- 111
        57488 => X"63",  -- 99
        57489 => X"54",  -- 84
        57490 => X"4B",  -- 75
        57491 => X"45",  -- 69
        57492 => X"40",  -- 64
        57493 => X"43",  -- 67
        57494 => X"61",  -- 97
        57495 => X"8B",  -- 139
        57496 => X"94",  -- 148
        57497 => X"90",  -- 144
        57498 => X"8E",  -- 142
        57499 => X"8E",  -- 142
        57500 => X"8E",  -- 142
        57501 => X"8E",  -- 142
        57502 => X"91",  -- 145
        57503 => X"95",  -- 149
        57504 => X"AC",  -- 172
        57505 => X"B5",  -- 181
        57506 => X"BB",  -- 187
        57507 => X"BA",  -- 186
        57508 => X"B7",  -- 183
        57509 => X"B9",  -- 185
        57510 => X"B9",  -- 185
        57511 => X"B8",  -- 184
        57512 => X"B0",  -- 176
        57513 => X"AB",  -- 171
        57514 => X"AA",  -- 170
        57515 => X"A4",  -- 164
        57516 => X"98",  -- 152
        57517 => X"99",  -- 153
        57518 => X"98",  -- 152
        57519 => X"91",  -- 145
        57520 => X"99",  -- 153
        57521 => X"B5",  -- 181
        57522 => X"B9",  -- 185
        57523 => X"C2",  -- 194
        57524 => X"99",  -- 153
        57525 => X"9A",  -- 154
        57526 => X"84",  -- 132
        57527 => X"82",  -- 130
        57528 => X"81",  -- 129
        57529 => X"8E",  -- 142
        57530 => X"A4",  -- 164
        57531 => X"A4",  -- 164
        57532 => X"B8",  -- 184
        57533 => X"BE",  -- 190
        57534 => X"CF",  -- 207
        57535 => X"CC",  -- 204
        57536 => X"BE",  -- 190
        57537 => X"BD",  -- 189
        57538 => X"AF",  -- 175
        57539 => X"9D",  -- 157
        57540 => X"A0",  -- 160
        57541 => X"9F",  -- 159
        57542 => X"95",  -- 149
        57543 => X"A0",  -- 160
        57544 => X"A3",  -- 163
        57545 => X"A6",  -- 166
        57546 => X"AD",  -- 173
        57547 => X"B7",  -- 183
        57548 => X"BD",  -- 189
        57549 => X"C1",  -- 193
        57550 => X"BE",  -- 190
        57551 => X"BB",  -- 187
        57552 => X"CA",  -- 202
        57553 => X"C0",  -- 192
        57554 => X"6E",  -- 110
        57555 => X"56",  -- 86
        57556 => X"62",  -- 98
        57557 => X"5E",  -- 94
        57558 => X"76",  -- 118
        57559 => X"74",  -- 116
        57560 => X"4D",  -- 77
        57561 => X"48",  -- 72
        57562 => X"59",  -- 89
        57563 => X"6A",  -- 106
        57564 => X"63",  -- 99
        57565 => X"59",  -- 89
        57566 => X"4D",  -- 77
        57567 => X"38",  -- 56
        57568 => X"30",  -- 48
        57569 => X"30",  -- 48
        57570 => X"2D",  -- 45
        57571 => X"33",  -- 51
        57572 => X"3D",  -- 61
        57573 => X"37",  -- 55
        57574 => X"2B",  -- 43
        57575 => X"2A",  -- 42
        57576 => X"2D",  -- 45
        57577 => X"2A",  -- 42
        57578 => X"2C",  -- 44
        57579 => X"33",  -- 51
        57580 => X"35",  -- 53
        57581 => X"37",  -- 55
        57582 => X"41",  -- 65
        57583 => X"4E",  -- 78
        57584 => X"44",  -- 68
        57585 => X"4D",  -- 77
        57586 => X"50",  -- 80
        57587 => X"4F",  -- 79
        57588 => X"5C",  -- 92
        57589 => X"6A",  -- 106
        57590 => X"61",  -- 97
        57591 => X"4A",  -- 74
        57592 => X"3B",  -- 59
        57593 => X"4F",  -- 79
        57594 => X"58",  -- 88
        57595 => X"57",  -- 87
        57596 => X"59",  -- 89
        57597 => X"5C",  -- 92
        57598 => X"64",  -- 100
        57599 => X"70",  -- 112
        57600 => X"27",  -- 39
        57601 => X"28",  -- 40
        57602 => X"27",  -- 39
        57603 => X"23",  -- 35
        57604 => X"22",  -- 34
        57605 => X"24",  -- 36
        57606 => X"23",  -- 35
        57607 => X"1F",  -- 31
        57608 => X"20",  -- 32
        57609 => X"1C",  -- 28
        57610 => X"1E",  -- 30
        57611 => X"24",  -- 36
        57612 => X"25",  -- 37
        57613 => X"23",  -- 35
        57614 => X"28",  -- 40
        57615 => X"33",  -- 51
        57616 => X"40",  -- 64
        57617 => X"42",  -- 66
        57618 => X"3B",  -- 59
        57619 => X"34",  -- 52
        57620 => X"30",  -- 48
        57621 => X"30",  -- 48
        57622 => X"2B",  -- 43
        57623 => X"23",  -- 35
        57624 => X"1D",  -- 29
        57625 => X"1C",  -- 28
        57626 => X"1B",  -- 27
        57627 => X"1C",  -- 28
        57628 => X"1D",  -- 29
        57629 => X"20",  -- 32
        57630 => X"23",  -- 35
        57631 => X"22",  -- 34
        57632 => X"27",  -- 39
        57633 => X"05",  -- 5
        57634 => X"23",  -- 35
        57635 => X"32",  -- 50
        57636 => X"21",  -- 33
        57637 => X"23",  -- 35
        57638 => X"26",  -- 38
        57639 => X"62",  -- 98
        57640 => X"AB",  -- 171
        57641 => X"84",  -- 132
        57642 => X"4D",  -- 77
        57643 => X"7B",  -- 123
        57644 => X"46",  -- 70
        57645 => X"38",  -- 56
        57646 => X"33",  -- 51
        57647 => X"43",  -- 67
        57648 => X"7A",  -- 122
        57649 => X"58",  -- 88
        57650 => X"3A",  -- 58
        57651 => X"43",  -- 67
        57652 => X"51",  -- 81
        57653 => X"4A",  -- 74
        57654 => X"75",  -- 117
        57655 => X"5F",  -- 95
        57656 => X"34",  -- 52
        57657 => X"37",  -- 55
        57658 => X"47",  -- 71
        57659 => X"6A",  -- 106
        57660 => X"77",  -- 119
        57661 => X"5B",  -- 91
        57662 => X"34",  -- 52
        57663 => X"27",  -- 39
        57664 => X"38",  -- 56
        57665 => X"50",  -- 80
        57666 => X"6E",  -- 110
        57667 => X"82",  -- 130
        57668 => X"7E",  -- 126
        57669 => X"63",  -- 99
        57670 => X"52",  -- 82
        57671 => X"59",  -- 89
        57672 => X"68",  -- 104
        57673 => X"5D",  -- 93
        57674 => X"5B",  -- 91
        57675 => X"6D",  -- 109
        57676 => X"86",  -- 134
        57677 => X"94",  -- 148
        57678 => X"95",  -- 149
        57679 => X"93",  -- 147
        57680 => X"8B",  -- 139
        57681 => X"86",  -- 134
        57682 => X"7C",  -- 124
        57683 => X"70",  -- 112
        57684 => X"5B",  -- 91
        57685 => X"3C",  -- 60
        57686 => X"18",  -- 24
        57687 => X"02",  -- 2
        57688 => X"15",  -- 21
        57689 => X"17",  -- 23
        57690 => X"1D",  -- 29
        57691 => X"20",  -- 32
        57692 => X"20",  -- 32
        57693 => X"1F",  -- 31
        57694 => X"1E",  -- 30
        57695 => X"21",  -- 33
        57696 => X"22",  -- 34
        57697 => X"1A",  -- 26
        57698 => X"10",  -- 16
        57699 => X"18",  -- 24
        57700 => X"3D",  -- 61
        57701 => X"6C",  -- 108
        57702 => X"86",  -- 134
        57703 => X"8B",  -- 139
        57704 => X"A4",  -- 164
        57705 => X"B2",  -- 178
        57706 => X"B5",  -- 181
        57707 => X"BF",  -- 191
        57708 => X"C3",  -- 195
        57709 => X"BF",  -- 191
        57710 => X"C2",  -- 194
        57711 => X"B5",  -- 181
        57712 => X"AB",  -- 171
        57713 => X"AA",  -- 170
        57714 => X"A7",  -- 167
        57715 => X"A7",  -- 167
        57716 => X"AD",  -- 173
        57717 => X"BC",  -- 188
        57718 => X"BB",  -- 187
        57719 => X"A4",  -- 164
        57720 => X"B1",  -- 177
        57721 => X"CB",  -- 203
        57722 => X"9D",  -- 157
        57723 => X"41",  -- 65
        57724 => X"4C",  -- 76
        57725 => X"83",  -- 131
        57726 => X"99",  -- 153
        57727 => X"C6",  -- 198
        57728 => X"99",  -- 153
        57729 => X"6A",  -- 106
        57730 => X"58",  -- 88
        57731 => X"47",  -- 71
        57732 => X"3D",  -- 61
        57733 => X"61",  -- 97
        57734 => X"88",  -- 136
        57735 => X"9E",  -- 158
        57736 => X"6B",  -- 107
        57737 => X"40",  -- 64
        57738 => X"34",  -- 52
        57739 => X"2D",  -- 45
        57740 => X"1B",  -- 27
        57741 => X"39",  -- 57
        57742 => X"2E",  -- 46
        57743 => X"19",  -- 25
        57744 => X"5E",  -- 94
        57745 => X"43",  -- 67
        57746 => X"23",  -- 35
        57747 => X"21",  -- 33
        57748 => X"19",  -- 25
        57749 => X"4F",  -- 79
        57750 => X"8C",  -- 140
        57751 => X"7D",  -- 125
        57752 => X"92",  -- 146
        57753 => X"72",  -- 114
        57754 => X"4F",  -- 79
        57755 => X"3D",  -- 61
        57756 => X"44",  -- 68
        57757 => X"51",  -- 81
        57758 => X"4F",  -- 79
        57759 => X"47",  -- 71
        57760 => X"49",  -- 73
        57761 => X"4B",  -- 75
        57762 => X"41",  -- 65
        57763 => X"36",  -- 54
        57764 => X"2A",  -- 42
        57765 => X"1D",  -- 29
        57766 => X"32",  -- 50
        57767 => X"62",  -- 98
        57768 => X"31",  -- 49
        57769 => X"1D",  -- 29
        57770 => X"24",  -- 36
        57771 => X"2E",  -- 46
        57772 => X"33",  -- 51
        57773 => X"3E",  -- 62
        57774 => X"39",  -- 57
        57775 => X"36",  -- 54
        57776 => X"32",  -- 50
        57777 => X"42",  -- 66
        57778 => X"63",  -- 99
        57779 => X"84",  -- 132
        57780 => X"88",  -- 136
        57781 => X"6E",  -- 110
        57782 => X"52",  -- 82
        57783 => X"45",  -- 69
        57784 => X"47",  -- 71
        57785 => X"3F",  -- 63
        57786 => X"32",  -- 50
        57787 => X"28",  -- 40
        57788 => X"22",  -- 34
        57789 => X"21",  -- 33
        57790 => X"26",  -- 38
        57791 => X"29",  -- 41
        57792 => X"2C",  -- 44
        57793 => X"38",  -- 56
        57794 => X"4D",  -- 77
        57795 => X"5F",  -- 95
        57796 => X"6B",  -- 107
        57797 => X"70",  -- 112
        57798 => X"70",  -- 112
        57799 => X"70",  -- 112
        57800 => X"76",  -- 118
        57801 => X"75",  -- 117
        57802 => X"72",  -- 114
        57803 => X"6E",  -- 110
        57804 => X"6C",  -- 108
        57805 => X"66",  -- 102
        57806 => X"60",  -- 96
        57807 => X"5D",  -- 93
        57808 => X"51",  -- 81
        57809 => X"41",  -- 65
        57810 => X"35",  -- 53
        57811 => X"33",  -- 51
        57812 => X"31",  -- 49
        57813 => X"41",  -- 65
        57814 => X"6B",  -- 107
        57815 => X"92",  -- 146
        57816 => X"8F",  -- 143
        57817 => X"8A",  -- 138
        57818 => X"8C",  -- 140
        57819 => X"98",  -- 152
        57820 => X"A0",  -- 160
        57821 => X"9E",  -- 158
        57822 => X"97",  -- 151
        57823 => X"91",  -- 145
        57824 => X"B9",  -- 185
        57825 => X"BA",  -- 186
        57826 => X"B9",  -- 185
        57827 => X"B6",  -- 182
        57828 => X"B4",  -- 180
        57829 => X"B3",  -- 179
        57830 => X"AF",  -- 175
        57831 => X"A9",  -- 169
        57832 => X"A9",  -- 169
        57833 => X"AA",  -- 170
        57834 => X"AE",  -- 174
        57835 => X"A9",  -- 169
        57836 => X"99",  -- 153
        57837 => X"94",  -- 148
        57838 => X"93",  -- 147
        57839 => X"8D",  -- 141
        57840 => X"94",  -- 148
        57841 => X"B1",  -- 177
        57842 => X"AC",  -- 172
        57843 => X"B0",  -- 176
        57844 => X"89",  -- 137
        57845 => X"8C",  -- 140
        57846 => X"7F",  -- 127
        57847 => X"8B",  -- 139
        57848 => X"8A",  -- 138
        57849 => X"94",  -- 148
        57850 => X"A4",  -- 164
        57851 => X"9A",  -- 154
        57852 => X"A5",  -- 165
        57853 => X"AB",  -- 171
        57854 => X"C0",  -- 192
        57855 => X"C3",  -- 195
        57856 => X"C8",  -- 200
        57857 => X"C8",  -- 200
        57858 => X"AF",  -- 175
        57859 => X"7E",  -- 126
        57860 => X"7A",  -- 122
        57861 => X"90",  -- 144
        57862 => X"93",  -- 147
        57863 => X"A1",  -- 161
        57864 => X"A0",  -- 160
        57865 => X"A2",  -- 162
        57866 => X"A7",  -- 167
        57867 => X"B1",  -- 177
        57868 => X"BA",  -- 186
        57869 => X"BF",  -- 191
        57870 => X"BF",  -- 191
        57871 => X"BE",  -- 190
        57872 => X"BC",  -- 188
        57873 => X"C4",  -- 196
        57874 => X"6D",  -- 109
        57875 => X"49",  -- 73
        57876 => X"5F",  -- 95
        57877 => X"4F",  -- 79
        57878 => X"52",  -- 82
        57879 => X"69",  -- 105
        57880 => X"5B",  -- 91
        57881 => X"43",  -- 67
        57882 => X"49",  -- 73
        57883 => X"5E",  -- 94
        57884 => X"59",  -- 89
        57885 => X"48",  -- 72
        57886 => X"3C",  -- 60
        57887 => X"2F",  -- 47
        57888 => X"2B",  -- 43
        57889 => X"2A",  -- 42
        57890 => X"25",  -- 37
        57891 => X"2A",  -- 42
        57892 => X"37",  -- 55
        57893 => X"35",  -- 53
        57894 => X"2B",  -- 43
        57895 => X"29",  -- 41
        57896 => X"27",  -- 39
        57897 => X"24",  -- 36
        57898 => X"28",  -- 40
        57899 => X"31",  -- 49
        57900 => X"35",  -- 53
        57901 => X"37",  -- 55
        57902 => X"3F",  -- 63
        57903 => X"4B",  -- 75
        57904 => X"4D",  -- 77
        57905 => X"5A",  -- 90
        57906 => X"58",  -- 88
        57907 => X"4A",  -- 74
        57908 => X"4C",  -- 76
        57909 => X"5D",  -- 93
        57910 => X"61",  -- 97
        57911 => X"57",  -- 87
        57912 => X"4C",  -- 76
        57913 => X"4D",  -- 77
        57914 => X"4F",  -- 79
        57915 => X"57",  -- 87
        57916 => X"5E",  -- 94
        57917 => X"5B",  -- 91
        57918 => X"64",  -- 100
        57919 => X"7B",  -- 123
        57920 => X"24",  -- 36
        57921 => X"25",  -- 37
        57922 => X"25",  -- 37
        57923 => X"22",  -- 34
        57924 => X"21",  -- 33
        57925 => X"23",  -- 35
        57926 => X"23",  -- 35
        57927 => X"1F",  -- 31
        57928 => X"24",  -- 36
        57929 => X"21",  -- 33
        57930 => X"22",  -- 34
        57931 => X"25",  -- 37
        57932 => X"28",  -- 40
        57933 => X"28",  -- 40
        57934 => X"29",  -- 41
        57935 => X"2B",  -- 43
        57936 => X"2F",  -- 47
        57937 => X"2D",  -- 45
        57938 => X"2B",  -- 43
        57939 => X"28",  -- 40
        57940 => X"2A",  -- 42
        57941 => X"2E",  -- 46
        57942 => X"2B",  -- 43
        57943 => X"24",  -- 36
        57944 => X"26",  -- 38
        57945 => X"23",  -- 35
        57946 => X"20",  -- 32
        57947 => X"1B",  -- 27
        57948 => X"19",  -- 25
        57949 => X"1A",  -- 26
        57950 => X"1C",  -- 28
        57951 => X"1D",  -- 29
        57952 => X"1C",  -- 28
        57953 => X"2D",  -- 45
        57954 => X"26",  -- 38
        57955 => X"0F",  -- 15
        57956 => X"2E",  -- 46
        57957 => X"47",  -- 71
        57958 => X"A0",  -- 160
        57959 => X"83",  -- 131
        57960 => X"30",  -- 48
        57961 => X"54",  -- 84
        57962 => X"6A",  -- 106
        57963 => X"39",  -- 57
        57964 => X"31",  -- 49
        57965 => X"48",  -- 72
        57966 => X"4A",  -- 74
        57967 => X"87",  -- 135
        57968 => X"58",  -- 88
        57969 => X"29",  -- 41
        57970 => X"57",  -- 87
        57971 => X"58",  -- 88
        57972 => X"62",  -- 98
        57973 => X"6D",  -- 109
        57974 => X"5E",  -- 94
        57975 => X"29",  -- 41
        57976 => X"41",  -- 65
        57977 => X"52",  -- 82
        57978 => X"5B",  -- 91
        57979 => X"57",  -- 87
        57980 => X"65",  -- 101
        57981 => X"63",  -- 99
        57982 => X"4F",  -- 79
        57983 => X"35",  -- 53
        57984 => X"2B",  -- 43
        57985 => X"27",  -- 39
        57986 => X"30",  -- 48
        57987 => X"4A",  -- 74
        57988 => X"56",  -- 86
        57989 => X"43",  -- 67
        57990 => X"37",  -- 55
        57991 => X"45",  -- 69
        57992 => X"67",  -- 103
        57993 => X"52",  -- 82
        57994 => X"38",  -- 56
        57995 => X"4C",  -- 76
        57996 => X"82",  -- 130
        57997 => X"9B",  -- 155
        57998 => X"95",  -- 149
        57999 => X"98",  -- 152
        58000 => X"93",  -- 147
        58001 => X"92",  -- 146
        58002 => X"89",  -- 137
        58003 => X"7A",  -- 122
        58004 => X"6F",  -- 111
        58005 => X"5B",  -- 91
        58006 => X"32",  -- 50
        58007 => X"0A",  -- 10
        58008 => X"14",  -- 20
        58009 => X"23",  -- 35
        58010 => X"28",  -- 40
        58011 => X"1B",  -- 27
        58012 => X"17",  -- 23
        58013 => X"1F",  -- 31
        58014 => X"22",  -- 34
        58015 => X"1C",  -- 28
        58016 => X"32",  -- 50
        58017 => X"10",  -- 16
        58018 => X"0F",  -- 15
        58019 => X"43",  -- 67
        58020 => X"7A",  -- 122
        58021 => X"8D",  -- 141
        58022 => X"94",  -- 148
        58023 => X"A1",  -- 161
        58024 => X"AD",  -- 173
        58025 => X"BF",  -- 191
        58026 => X"C2",  -- 194
        58027 => X"C5",  -- 197
        58028 => X"BE",  -- 190
        58029 => X"B6",  -- 182
        58030 => X"BA",  -- 186
        58031 => X"B2",  -- 178
        58032 => X"A2",  -- 162
        58033 => X"97",  -- 151
        58034 => X"7A",  -- 122
        58035 => X"8D",  -- 141
        58036 => X"A5",  -- 165
        58037 => X"AC",  -- 172
        58038 => X"AF",  -- 175
        58039 => X"83",  -- 131
        58040 => X"63",  -- 99
        58041 => X"5F",  -- 95
        58042 => X"56",  -- 86
        58043 => X"69",  -- 105
        58044 => X"A0",  -- 160
        58045 => X"AE",  -- 174
        58046 => X"97",  -- 151
        58047 => X"A2",  -- 162
        58048 => X"8A",  -- 138
        58049 => X"54",  -- 84
        58050 => X"49",  -- 73
        58051 => X"3D",  -- 61
        58052 => X"37",  -- 55
        58053 => X"3F",  -- 63
        58054 => X"35",  -- 53
        58055 => X"3C",  -- 60
        58056 => X"7A",  -- 122
        58057 => X"8A",  -- 138
        58058 => X"6A",  -- 106
        58059 => X"4C",  -- 76
        58060 => X"1D",  -- 29
        58061 => X"29",  -- 41
        58062 => X"3F",  -- 63
        58063 => X"1E",  -- 30
        58064 => X"1B",  -- 27
        58065 => X"61",  -- 97
        58066 => X"44",  -- 68
        58067 => X"0E",  -- 14
        58068 => X"20",  -- 32
        58069 => X"2C",  -- 44
        58070 => X"37",  -- 55
        58071 => X"59",  -- 89
        58072 => X"77",  -- 119
        58073 => X"8B",  -- 139
        58074 => X"8E",  -- 142
        58075 => X"5F",  -- 95
        58076 => X"3A",  -- 58
        58077 => X"3D",  -- 61
        58078 => X"42",  -- 66
        58079 => X"4B",  -- 75
        58080 => X"50",  -- 80
        58081 => X"47",  -- 71
        58082 => X"3E",  -- 62
        58083 => X"3C",  -- 60
        58084 => X"37",  -- 55
        58085 => X"26",  -- 38
        58086 => X"26",  -- 38
        58087 => X"39",  -- 57
        58088 => X"81",  -- 129
        58089 => X"33",  -- 51
        58090 => X"28",  -- 40
        58091 => X"37",  -- 55
        58092 => X"30",  -- 48
        58093 => X"33",  -- 51
        58094 => X"34",  -- 52
        58095 => X"29",  -- 41
        58096 => X"31",  -- 49
        58097 => X"2C",  -- 44
        58098 => X"2D",  -- 45
        58099 => X"3A",  -- 58
        58100 => X"4C",  -- 76
        58101 => X"61",  -- 97
        58102 => X"7B",  -- 123
        58103 => X"90",  -- 144
        58104 => X"6E",  -- 110
        58105 => X"63",  -- 99
        58106 => X"54",  -- 84
        58107 => X"4B",  -- 75
        58108 => X"47",  -- 71
        58109 => X"47",  -- 71
        58110 => X"4E",  -- 78
        58111 => X"54",  -- 84
        58112 => X"6D",  -- 109
        58113 => X"63",  -- 99
        58114 => X"59",  -- 89
        58115 => X"5A",  -- 90
        58116 => X"5F",  -- 95
        58117 => X"64",  -- 100
        58118 => X"67",  -- 103
        58119 => X"68",  -- 104
        58120 => X"6F",  -- 111
        58121 => X"6C",  -- 108
        58122 => X"67",  -- 103
        58123 => X"60",  -- 96
        58124 => X"5A",  -- 90
        58125 => X"53",  -- 83
        58126 => X"4A",  -- 74
        58127 => X"46",  -- 70
        58128 => X"45",  -- 69
        58129 => X"3A",  -- 58
        58130 => X"2C",  -- 44
        58131 => X"2E",  -- 46
        58132 => X"31",  -- 49
        58133 => X"47",  -- 71
        58134 => X"76",  -- 118
        58135 => X"8C",  -- 140
        58136 => X"88",  -- 136
        58137 => X"8E",  -- 142
        58138 => X"94",  -- 148
        58139 => X"96",  -- 150
        58140 => X"93",  -- 147
        58141 => X"92",  -- 146
        58142 => X"99",  -- 153
        58143 => X"A3",  -- 163
        58144 => X"B1",  -- 177
        58145 => X"AF",  -- 175
        58146 => X"AB",  -- 171
        58147 => X"A5",  -- 165
        58148 => X"9F",  -- 159
        58149 => X"98",  -- 152
        58150 => X"92",  -- 146
        58151 => X"8E",  -- 142
        58152 => X"8E",  -- 142
        58153 => X"97",  -- 151
        58154 => X"A8",  -- 168
        58155 => X"AA",  -- 170
        58156 => X"9E",  -- 158
        58157 => X"98",  -- 152
        58158 => X"90",  -- 144
        58159 => X"84",  -- 132
        58160 => X"A4",  -- 164
        58161 => X"A9",  -- 169
        58162 => X"90",  -- 144
        58163 => X"8A",  -- 138
        58164 => X"7F",  -- 127
        58165 => X"92",  -- 146
        58166 => X"91",  -- 145
        58167 => X"A3",  -- 163
        58168 => X"91",  -- 145
        58169 => X"9C",  -- 156
        58170 => X"AA",  -- 170
        58171 => X"AC",  -- 172
        58172 => X"B2",  -- 178
        58173 => X"AF",  -- 175
        58174 => X"B3",  -- 179
        58175 => X"B1",  -- 177
        58176 => X"C3",  -- 195
        58177 => X"D0",  -- 208
        58178 => X"C3",  -- 195
        58179 => X"7D",  -- 125
        58180 => X"64",  -- 100
        58181 => X"87",  -- 135
        58182 => X"9D",  -- 157
        58183 => X"B8",  -- 184
        58184 => X"B4",  -- 180
        58185 => X"B0",  -- 176
        58186 => X"AD",  -- 173
        58187 => X"AF",  -- 175
        58188 => X"B5",  -- 181
        58189 => X"BC",  -- 188
        58190 => X"C1",  -- 193
        58191 => X"C2",  -- 194
        58192 => X"C2",  -- 194
        58193 => X"C5",  -- 197
        58194 => X"6B",  -- 107
        58195 => X"33",  -- 51
        58196 => X"50",  -- 80
        58197 => X"50",  -- 80
        58198 => X"46",  -- 70
        58199 => X"61",  -- 97
        58200 => X"52",  -- 82
        58201 => X"3C",  -- 60
        58202 => X"3A",  -- 58
        58203 => X"4F",  -- 79
        58204 => X"51",  -- 81
        58205 => X"3F",  -- 63
        58206 => X"30",  -- 48
        58207 => X"29",  -- 41
        58208 => X"2A",  -- 42
        58209 => X"29",  -- 41
        58210 => X"23",  -- 35
        58211 => X"25",  -- 37
        58212 => X"30",  -- 48
        58213 => X"30",  -- 48
        58214 => X"28",  -- 40
        58215 => X"27",  -- 39
        58216 => X"1D",  -- 29
        58217 => X"1E",  -- 30
        58218 => X"24",  -- 36
        58219 => X"2D",  -- 45
        58220 => X"34",  -- 52
        58221 => X"38",  -- 56
        58222 => X"3C",  -- 60
        58223 => X"41",  -- 65
        58224 => X"45",  -- 69
        58225 => X"56",  -- 86
        58226 => X"59",  -- 89
        58227 => X"4D",  -- 77
        58228 => X"45",  -- 69
        58229 => X"4E",  -- 78
        58230 => X"59",  -- 89
        58231 => X"5C",  -- 92
        58232 => X"5D",  -- 93
        58233 => X"53",  -- 83
        58234 => X"4E",  -- 78
        58235 => X"5A",  -- 90
        58236 => X"64",  -- 100
        58237 => X"5F",  -- 95
        58238 => X"68",  -- 104
        58239 => X"82",  -- 130
        58240 => X"21",  -- 33
        58241 => X"23",  -- 35
        58242 => X"24",  -- 36
        58243 => X"22",  -- 34
        58244 => X"23",  -- 35
        58245 => X"27",  -- 39
        58246 => X"27",  -- 39
        58247 => X"24",  -- 36
        58248 => X"27",  -- 39
        58249 => X"29",  -- 41
        58250 => X"2A",  -- 42
        58251 => X"28",  -- 40
        58252 => X"26",  -- 38
        58253 => X"28",  -- 40
        58254 => X"26",  -- 38
        58255 => X"24",  -- 36
        58256 => X"1E",  -- 30
        58257 => X"1D",  -- 29
        58258 => X"1C",  -- 28
        58259 => X"1E",  -- 30
        58260 => X"26",  -- 38
        58261 => X"2E",  -- 46
        58262 => X"2C",  -- 44
        58263 => X"26",  -- 38
        58264 => X"2E",  -- 46
        58265 => X"2A",  -- 42
        58266 => X"24",  -- 36
        58267 => X"1C",  -- 28
        58268 => X"19",  -- 25
        58269 => X"17",  -- 23
        58270 => X"1A",  -- 26
        58271 => X"1C",  -- 28
        58272 => X"1F",  -- 31
        58273 => X"1F",  -- 31
        58274 => X"21",  -- 33
        58275 => X"6A",  -- 106
        58276 => X"90",  -- 144
        58277 => X"63",  -- 99
        58278 => X"77",  -- 119
        58279 => X"35",  -- 53
        58280 => X"83",  -- 131
        58281 => X"43",  -- 67
        58282 => X"31",  -- 49
        58283 => X"30",  -- 48
        58284 => X"29",  -- 41
        58285 => X"53",  -- 83
        58286 => X"80",  -- 128
        58287 => X"3C",  -- 60
        58288 => X"54",  -- 84
        58289 => X"80",  -- 128
        58290 => X"85",  -- 133
        58291 => X"79",  -- 121
        58292 => X"87",  -- 135
        58293 => X"39",  -- 57
        58294 => X"39",  -- 57
        58295 => X"60",  -- 96
        58296 => X"5B",  -- 91
        58297 => X"49",  -- 73
        58298 => X"37",  -- 55
        58299 => X"2B",  -- 43
        58300 => X"6A",  -- 106
        58301 => X"8C",  -- 140
        58302 => X"8A",  -- 138
        58303 => X"67",  -- 103
        58304 => X"55",  -- 85
        58305 => X"37",  -- 55
        58306 => X"1E",  -- 30
        58307 => X"24",  -- 36
        58308 => X"30",  -- 48
        58309 => X"2B",  -- 43
        58310 => X"30",  -- 48
        58311 => X"49",  -- 73
        58312 => X"71",  -- 113
        58313 => X"5E",  -- 94
        58314 => X"4D",  -- 77
        58315 => X"5D",  -- 93
        58316 => X"83",  -- 131
        58317 => X"91",  -- 145
        58318 => X"8C",  -- 140
        58319 => X"8B",  -- 139
        58320 => X"98",  -- 152
        58321 => X"99",  -- 153
        58322 => X"91",  -- 145
        58323 => X"85",  -- 133
        58324 => X"7F",  -- 127
        58325 => X"74",  -- 116
        58326 => X"53",  -- 83
        58327 => X"31",  -- 49
        58328 => X"19",  -- 25
        58329 => X"25",  -- 37
        58330 => X"29",  -- 41
        58331 => X"1D",  -- 29
        58332 => X"16",  -- 22
        58333 => X"1D",  -- 29
        58334 => X"26",  -- 38
        58335 => X"28",  -- 40
        58336 => X"3B",  -- 59
        58337 => X"1E",  -- 30
        58338 => X"2B",  -- 43
        58339 => X"6D",  -- 109
        58340 => X"A2",  -- 162
        58341 => X"A5",  -- 165
        58342 => X"A2",  -- 162
        58343 => X"AE",  -- 174
        58344 => X"BC",  -- 188
        58345 => X"BD",  -- 189
        58346 => X"B5",  -- 181
        58347 => X"B5",  -- 181
        58348 => X"A7",  -- 167
        58349 => X"9A",  -- 154
        58350 => X"B1",  -- 177
        58351 => X"C4",  -- 196
        58352 => X"A9",  -- 169
        58353 => X"7B",  -- 123
        58354 => X"48",  -- 72
        58355 => X"64",  -- 100
        58356 => X"8C",  -- 140
        58357 => X"92",  -- 146
        58358 => X"82",  -- 130
        58359 => X"4B",  -- 75
        58360 => X"2A",  -- 42
        58361 => X"47",  -- 71
        58362 => X"71",  -- 113
        58363 => X"A1",  -- 161
        58364 => X"B8",  -- 184
        58365 => X"C2",  -- 194
        58366 => X"C5",  -- 197
        58367 => X"B5",  -- 181
        58368 => X"71",  -- 113
        58369 => X"3E",  -- 62
        58370 => X"4A",  -- 74
        58371 => X"5B",  -- 91
        58372 => X"3D",  -- 61
        58373 => X"35",  -- 53
        58374 => X"47",  -- 71
        58375 => X"45",  -- 69
        58376 => X"1E",  -- 30
        58377 => X"20",  -- 32
        58378 => X"74",  -- 116
        58379 => X"86",  -- 134
        58380 => X"53",  -- 83
        58381 => X"43",  -- 67
        58382 => X"19",  -- 25
        58383 => X"34",  -- 52
        58384 => X"0C",  -- 12
        58385 => X"23",  -- 35
        58386 => X"51",  -- 81
        58387 => X"3B",  -- 59
        58388 => X"2E",  -- 46
        58389 => X"23",  -- 35
        58390 => X"36",  -- 54
        58391 => X"37",  -- 55
        58392 => X"3C",  -- 60
        58393 => X"4A",  -- 74
        58394 => X"82",  -- 130
        58395 => X"9B",  -- 155
        58396 => X"7B",  -- 123
        58397 => X"41",  -- 65
        58398 => X"22",  -- 34
        58399 => X"3F",  -- 63
        58400 => X"34",  -- 52
        58401 => X"41",  -- 65
        58402 => X"4B",  -- 75
        58403 => X"3A",  -- 58
        58404 => X"26",  -- 38
        58405 => X"32",  -- 50
        58406 => X"38",  -- 56
        58407 => X"23",  -- 35
        58408 => X"30",  -- 48
        58409 => X"68",  -- 104
        58410 => X"58",  -- 88
        58411 => X"26",  -- 38
        58412 => X"3A",  -- 58
        58413 => X"3F",  -- 63
        58414 => X"23",  -- 35
        58415 => X"39",  -- 57
        58416 => X"2C",  -- 44
        58417 => X"33",  -- 51
        58418 => X"3F",  -- 63
        58419 => X"4A",  -- 74
        58420 => X"52",  -- 82
        58421 => X"4F",  -- 79
        58422 => X"45",  -- 69
        58423 => X"3E",  -- 62
        58424 => X"61",  -- 97
        58425 => X"58",  -- 88
        58426 => X"50",  -- 80
        58427 => X"4A",  -- 74
        58428 => X"46",  -- 70
        58429 => X"48",  -- 72
        58430 => X"50",  -- 80
        58431 => X"5B",  -- 91
        58432 => X"46",  -- 70
        58433 => X"3E",  -- 62
        58434 => X"41",  -- 65
        58435 => X"57",  -- 87
        58436 => X"6E",  -- 110
        58437 => X"77",  -- 119
        58438 => X"74",  -- 116
        58439 => X"6E",  -- 110
        58440 => X"64",  -- 100
        58441 => X"60",  -- 96
        58442 => X"59",  -- 89
        58443 => X"51",  -- 81
        58444 => X"4B",  -- 75
        58445 => X"45",  -- 69
        58446 => X"3F",  -- 63
        58447 => X"3A",  -- 58
        58448 => X"3D",  -- 61
        58449 => X"38",  -- 56
        58450 => X"2B",  -- 43
        58451 => X"31",  -- 49
        58452 => X"38",  -- 56
        58453 => X"51",  -- 81
        58454 => X"7D",  -- 125
        58455 => X"7E",  -- 126
        58456 => X"86",  -- 134
        58457 => X"92",  -- 146
        58458 => X"98",  -- 152
        58459 => X"8A",  -- 138
        58460 => X"7B",  -- 123
        58461 => X"82",  -- 130
        58462 => X"9F",  -- 159
        58463 => X"B9",  -- 185
        58464 => X"A7",  -- 167
        58465 => X"A2",  -- 162
        58466 => X"97",  -- 151
        58467 => X"89",  -- 137
        58468 => X"7B",  -- 123
        58469 => X"75",  -- 117
        58470 => X"77",  -- 119
        58471 => X"7C",  -- 124
        58472 => X"85",  -- 133
        58473 => X"8F",  -- 143
        58474 => X"A1",  -- 161
        58475 => X"AC",  -- 172
        58476 => X"A6",  -- 166
        58477 => X"9E",  -- 158
        58478 => X"8E",  -- 142
        58479 => X"7C",  -- 124
        58480 => X"97",  -- 151
        58481 => X"9A",  -- 154
        58482 => X"8D",  -- 141
        58483 => X"92",  -- 146
        58484 => X"A2",  -- 162
        58485 => X"A8",  -- 168
        58486 => X"97",  -- 151
        58487 => X"92",  -- 146
        58488 => X"90",  -- 144
        58489 => X"94",  -- 148
        58490 => X"9F",  -- 159
        58491 => X"B3",  -- 179
        58492 => X"BB",  -- 187
        58493 => X"BC",  -- 188
        58494 => X"AE",  -- 174
        58495 => X"A8",  -- 168
        58496 => X"BB",  -- 187
        58497 => X"CE",  -- 206
        58498 => X"D8",  -- 216
        58499 => X"90",  -- 144
        58500 => X"65",  -- 101
        58501 => X"8A",  -- 138
        58502 => X"A8",  -- 168
        58503 => X"C4",  -- 196
        58504 => X"C3",  -- 195
        58505 => X"BF",  -- 191
        58506 => X"BB",  -- 187
        58507 => X"B9",  -- 185
        58508 => X"BA",  -- 186
        58509 => X"BD",  -- 189
        58510 => X"C1",  -- 193
        58511 => X"C5",  -- 197
        58512 => X"CB",  -- 203
        58513 => X"C3",  -- 195
        58514 => X"7E",  -- 126
        58515 => X"2B",  -- 43
        58516 => X"30",  -- 48
        58517 => X"4F",  -- 79
        58518 => X"4B",  -- 75
        58519 => X"59",  -- 89
        58520 => X"42",  -- 66
        58521 => X"38",  -- 56
        58522 => X"2F",  -- 47
        58523 => X"37",  -- 55
        58524 => X"45",  -- 69
        58525 => X"40",  -- 64
        58526 => X"31",  -- 49
        58527 => X"2A",  -- 42
        58528 => X"26",  -- 38
        58529 => X"29",  -- 41
        58530 => X"24",  -- 36
        58531 => X"23",  -- 35
        58532 => X"2A",  -- 42
        58533 => X"29",  -- 41
        58534 => X"23",  -- 35
        58535 => X"24",  -- 36
        58536 => X"1B",  -- 27
        58537 => X"1C",  -- 28
        58538 => X"1C",  -- 28
        58539 => X"20",  -- 32
        58540 => X"2A",  -- 42
        58541 => X"36",  -- 54
        58542 => X"3C",  -- 60
        58543 => X"3C",  -- 60
        58544 => X"37",  -- 55
        58545 => X"45",  -- 69
        58546 => X"51",  -- 81
        58547 => X"4F",  -- 79
        58548 => X"48",  -- 72
        58549 => X"48",  -- 72
        58550 => X"52",  -- 82
        58551 => X"5D",  -- 93
        58552 => X"61",  -- 97
        58553 => X"5B",  -- 91
        58554 => X"57",  -- 87
        58555 => X"60",  -- 96
        58556 => X"6A",  -- 106
        58557 => X"69",  -- 105
        58558 => X"71",  -- 113
        58559 => X"87",  -- 135
        58560 => X"20",  -- 32
        58561 => X"22",  -- 34
        58562 => X"23",  -- 35
        58563 => X"24",  -- 36
        58564 => X"27",  -- 39
        58565 => X"2C",  -- 44
        58566 => X"2D",  -- 45
        58567 => X"2A",  -- 42
        58568 => X"29",  -- 41
        58569 => X"2F",  -- 47
        58570 => X"30",  -- 48
        58571 => X"2A",  -- 42
        58572 => X"25",  -- 37
        58573 => X"25",  -- 37
        58574 => X"23",  -- 35
        58575 => X"1D",  -- 29
        58576 => X"1B",  -- 27
        58577 => X"19",  -- 25
        58578 => X"18",  -- 24
        58579 => X"1D",  -- 29
        58580 => X"26",  -- 38
        58581 => X"2E",  -- 46
        58582 => X"2D",  -- 45
        58583 => X"27",  -- 39
        58584 => X"30",  -- 48
        58585 => X"2C",  -- 44
        58586 => X"25",  -- 37
        58587 => X"1E",  -- 30
        58588 => X"1B",  -- 27
        58589 => X"1C",  -- 28
        58590 => X"1F",  -- 31
        58591 => X"22",  -- 34
        58592 => X"28",  -- 40
        58593 => X"4A",  -- 74
        58594 => X"88",  -- 136
        58595 => X"61",  -- 97
        58596 => X"1E",  -- 30
        58597 => X"66",  -- 102
        58598 => X"5A",  -- 90
        58599 => X"75",  -- 117
        58600 => X"31",  -- 49
        58601 => X"24",  -- 36
        58602 => X"28",  -- 40
        58603 => X"32",  -- 50
        58604 => X"5E",  -- 94
        58605 => X"7D",  -- 125
        58606 => X"5A",  -- 90
        58607 => X"99",  -- 153
        58608 => X"A0",  -- 160
        58609 => X"7B",  -- 123
        58610 => X"82",  -- 130
        58611 => X"57",  -- 87
        58612 => X"4F",  -- 79
        58613 => X"56",  -- 86
        58614 => X"6A",  -- 106
        58615 => X"3E",  -- 62
        58616 => X"35",  -- 53
        58617 => X"2D",  -- 45
        58618 => X"36",  -- 54
        58619 => X"30",  -- 48
        58620 => X"64",  -- 100
        58621 => X"6D",  -- 109
        58622 => X"7F",  -- 127
        58623 => X"79",  -- 121
        58624 => X"7A",  -- 122
        58625 => X"6D",  -- 109
        58626 => X"59",  -- 89
        58627 => X"43",  -- 67
        58628 => X"2D",  -- 45
        58629 => X"1A",  -- 26
        58630 => X"29",  -- 41
        58631 => X"4D",  -- 77
        58632 => X"4C",  -- 76
        58633 => X"53",  -- 83
        58634 => X"6A",  -- 106
        58635 => X"85",  -- 133
        58636 => X"92",  -- 146
        58637 => X"94",  -- 148
        58638 => X"95",  -- 149
        58639 => X"91",  -- 145
        58640 => X"9B",  -- 155
        58641 => X"9C",  -- 156
        58642 => X"97",  -- 151
        58643 => X"90",  -- 144
        58644 => X"8C",  -- 140
        58645 => X"86",  -- 134
        58646 => X"6F",  -- 111
        58647 => X"57",  -- 87
        58648 => X"1F",  -- 31
        58649 => X"1E",  -- 30
        58650 => X"21",  -- 33
        58651 => X"22",  -- 34
        58652 => X"17",  -- 23
        58653 => X"0E",  -- 14
        58654 => X"18",  -- 24
        58655 => X"2D",  -- 45
        58656 => X"23",  -- 35
        58657 => X"2E",  -- 46
        58658 => X"52",  -- 82
        58659 => X"82",  -- 130
        58660 => X"9B",  -- 155
        58661 => X"9F",  -- 159
        58662 => X"A8",  -- 168
        58663 => X"B9",  -- 185
        58664 => X"B3",  -- 179
        58665 => X"C2",  -- 194
        58666 => X"C3",  -- 195
        58667 => X"BB",  -- 187
        58668 => X"A3",  -- 163
        58669 => X"91",  -- 145
        58670 => X"9C",  -- 156
        58671 => X"A3",  -- 163
        58672 => X"90",  -- 144
        58673 => X"82",  -- 130
        58674 => X"6A",  -- 106
        58675 => X"59",  -- 89
        58676 => X"43",  -- 67
        58677 => X"3C",  -- 60
        58678 => X"4F",  -- 79
        58679 => X"51",  -- 81
        58680 => X"62",  -- 98
        58681 => X"92",  -- 146
        58682 => X"93",  -- 147
        58683 => X"A9",  -- 169
        58684 => X"CB",  -- 203
        58685 => X"B8",  -- 184
        58686 => X"9F",  -- 159
        58687 => X"8E",  -- 142
        58688 => X"AA",  -- 170
        58689 => X"BB",  -- 187
        58690 => X"8C",  -- 140
        58691 => X"60",  -- 96
        58692 => X"46",  -- 70
        58693 => X"29",  -- 41
        58694 => X"33",  -- 51
        58695 => X"47",  -- 71
        58696 => X"59",  -- 89
        58697 => X"52",  -- 82
        58698 => X"0D",  -- 13
        58699 => X"21",  -- 33
        58700 => X"82",  -- 130
        58701 => X"8C",  -- 140
        58702 => X"40",  -- 64
        58703 => X"46",  -- 70
        58704 => X"4B",  -- 75
        58705 => X"16",  -- 22
        58706 => X"35",  -- 53
        58707 => X"62",  -- 98
        58708 => X"20",  -- 32
        58709 => X"2E",  -- 46
        58710 => X"2F",  -- 47
        58711 => X"32",  -- 50
        58712 => X"3D",  -- 61
        58713 => X"33",  -- 51
        58714 => X"40",  -- 64
        58715 => X"51",  -- 81
        58716 => X"7E",  -- 126
        58717 => X"93",  -- 147
        58718 => X"58",  -- 88
        58719 => X"1E",  -- 30
        58720 => X"27",  -- 39
        58721 => X"2B",  -- 43
        58722 => X"2D",  -- 45
        58723 => X"34",  -- 52
        58724 => X"37",  -- 55
        58725 => X"2B",  -- 43
        58726 => X"23",  -- 35
        58727 => X"29",  -- 41
        58728 => X"23",  -- 35
        58729 => X"40",  -- 64
        58730 => X"73",  -- 115
        58731 => X"5E",  -- 94
        58732 => X"2B",  -- 43
        58733 => X"2B",  -- 43
        58734 => X"33",  -- 51
        58735 => X"27",  -- 39
        58736 => X"2C",  -- 44
        58737 => X"2E",  -- 46
        58738 => X"32",  -- 50
        58739 => X"3C",  -- 60
        58740 => X"4B",  -- 75
        58741 => X"57",  -- 87
        58742 => X"57",  -- 87
        58743 => X"50",  -- 80
        58744 => X"4E",  -- 78
        58745 => X"4C",  -- 76
        58746 => X"4A",  -- 74
        58747 => X"47",  -- 71
        58748 => X"43",  -- 67
        58749 => X"42",  -- 66
        58750 => X"4F",  -- 79
        58751 => X"5D",  -- 93
        58752 => X"65",  -- 101
        58753 => X"55",  -- 85
        58754 => X"4E",  -- 78
        58755 => X"5D",  -- 93
        58756 => X"74",  -- 116
        58757 => X"7B",  -- 123
        58758 => X"74",  -- 116
        58759 => X"6A",  -- 106
        58760 => X"5E",  -- 94
        58761 => X"59",  -- 89
        58762 => X"52",  -- 82
        58763 => X"4A",  -- 74
        58764 => X"46",  -- 70
        58765 => X"41",  -- 65
        58766 => X"3D",  -- 61
        58767 => X"3A",  -- 58
        58768 => X"35",  -- 53
        58769 => X"35",  -- 53
        58770 => X"2B",  -- 43
        58771 => X"34",  -- 52
        58772 => X"3C",  -- 60
        58773 => X"59",  -- 89
        58774 => X"7E",  -- 126
        58775 => X"73",  -- 115
        58776 => X"89",  -- 137
        58777 => X"92",  -- 146
        58778 => X"90",  -- 144
        58779 => X"86",  -- 134
        58780 => X"82",  -- 130
        58781 => X"90",  -- 144
        58782 => X"A7",  -- 167
        58783 => X"B5",  -- 181
        58784 => X"A5",  -- 165
        58785 => X"9D",  -- 157
        58786 => X"8B",  -- 139
        58787 => X"74",  -- 116
        58788 => X"60",  -- 96
        58789 => X"5F",  -- 95
        58790 => X"6F",  -- 111
        58791 => X"80",  -- 128
        58792 => X"98",  -- 152
        58793 => X"9B",  -- 155
        58794 => X"A9",  -- 169
        58795 => X"B1",  -- 177
        58796 => X"AF",  -- 175
        58797 => X"A7",  -- 167
        58798 => X"94",  -- 148
        58799 => X"7B",  -- 123
        58800 => X"8B",  -- 139
        58801 => X"9B",  -- 155
        58802 => X"9F",  -- 159
        58803 => X"A2",  -- 162
        58804 => X"B0",  -- 176
        58805 => X"AB",  -- 171
        58806 => X"9E",  -- 158
        58807 => X"9F",  -- 159
        58808 => X"A3",  -- 163
        58809 => X"98",  -- 152
        58810 => X"8B",  -- 139
        58811 => X"A4",  -- 164
        58812 => X"AC",  -- 172
        58813 => X"B8",  -- 184
        58814 => X"AB",  -- 171
        58815 => X"AB",  -- 171
        58816 => X"B1",  -- 177
        58817 => X"BF",  -- 191
        58818 => X"D7",  -- 215
        58819 => X"9B",  -- 155
        58820 => X"70",  -- 112
        58821 => X"95",  -- 149
        58822 => X"AF",  -- 175
        58823 => X"C3",  -- 195
        58824 => X"BF",  -- 191
        58825 => X"C0",  -- 192
        58826 => X"BF",  -- 191
        58827 => X"C0",  -- 192
        58828 => X"BF",  -- 191
        58829 => X"BE",  -- 190
        58830 => X"BE",  -- 190
        58831 => X"BF",  -- 191
        58832 => X"C8",  -- 200
        58833 => X"C2",  -- 194
        58834 => X"9C",  -- 156
        58835 => X"38",  -- 56
        58836 => X"1C",  -- 28
        58837 => X"49",  -- 73
        58838 => X"47",  -- 71
        58839 => X"40",  -- 64
        58840 => X"42",  -- 66
        58841 => X"40",  -- 64
        58842 => X"2C",  -- 44
        58843 => X"25",  -- 37
        58844 => X"37",  -- 55
        58845 => X"3D",  -- 61
        58846 => X"2F",  -- 47
        58847 => X"28",  -- 40
        58848 => X"23",  -- 35
        58849 => X"29",  -- 41
        58850 => X"25",  -- 37
        58851 => X"22",  -- 34
        58852 => X"26",  -- 38
        58853 => X"24",  -- 36
        58854 => X"1F",  -- 31
        58855 => X"20",  -- 32
        58856 => X"20",  -- 32
        58857 => X"1C",  -- 28
        58858 => X"14",  -- 20
        58859 => X"11",  -- 17
        58860 => X"1D",  -- 29
        58861 => X"32",  -- 50
        58862 => X"3E",  -- 62
        58863 => X"3E",  -- 62
        58864 => X"36",  -- 54
        58865 => X"3E",  -- 62
        58866 => X"4B",  -- 75
        58867 => X"51",  -- 81
        58868 => X"4B",  -- 75
        58869 => X"44",  -- 68
        58870 => X"4B",  -- 75
        58871 => X"59",  -- 89
        58872 => X"60",  -- 96
        58873 => X"63",  -- 99
        58874 => X"63",  -- 99
        58875 => X"68",  -- 104
        58876 => X"72",  -- 114
        58877 => X"75",  -- 117
        58878 => X"7C",  -- 124
        58879 => X"8C",  -- 140
        58880 => X"22",  -- 34
        58881 => X"26",  -- 38
        58882 => X"27",  -- 39
        58883 => X"26",  -- 38
        58884 => X"29",  -- 41
        58885 => X"2E",  -- 46
        58886 => X"31",  -- 49
        58887 => X"2F",  -- 47
        58888 => X"31",  -- 49
        58889 => X"2F",  -- 47
        58890 => X"2B",  -- 43
        58891 => X"25",  -- 37
        58892 => X"21",  -- 33
        58893 => X"1E",  -- 30
        58894 => X"1C",  -- 28
        58895 => X"1B",  -- 27
        58896 => X"22",  -- 34
        58897 => X"1C",  -- 28
        58898 => X"17",  -- 23
        58899 => X"1C",  -- 28
        58900 => X"27",  -- 39
        58901 => X"2E",  -- 46
        58902 => X"2A",  -- 42
        58903 => X"24",  -- 36
        58904 => X"2C",  -- 44
        58905 => X"3F",  -- 63
        58906 => X"29",  -- 41
        58907 => X"20",  -- 32
        58908 => X"2F",  -- 47
        58909 => X"27",  -- 39
        58910 => X"26",  -- 38
        58911 => X"3C",  -- 60
        58912 => X"6B",  -- 107
        58913 => X"84",  -- 132
        58914 => X"2B",  -- 43
        58915 => X"1E",  -- 30
        58916 => X"48",  -- 72
        58917 => X"80",  -- 128
        58918 => X"60",  -- 96
        58919 => X"29",  -- 41
        58920 => X"26",  -- 38
        58921 => X"2A",  -- 42
        58922 => X"2A",  -- 42
        58923 => X"4E",  -- 78
        58924 => X"7D",  -- 125
        58925 => X"98",  -- 152
        58926 => X"9C",  -- 156
        58927 => X"81",  -- 129
        58928 => X"67",  -- 103
        58929 => X"65",  -- 101
        58930 => X"48",  -- 72
        58931 => X"62",  -- 98
        58932 => X"70",  -- 112
        58933 => X"51",  -- 81
        58934 => X"2A",  -- 42
        58935 => X"37",  -- 55
        58936 => X"41",  -- 65
        58937 => X"6A",  -- 106
        58938 => X"29",  -- 41
        58939 => X"29",  -- 41
        58940 => X"4A",  -- 74
        58941 => X"44",  -- 68
        58942 => X"67",  -- 103
        58943 => X"88",  -- 136
        58944 => X"87",  -- 135
        58945 => X"7F",  -- 127
        58946 => X"84",  -- 132
        58947 => X"68",  -- 104
        58948 => X"55",  -- 85
        58949 => X"4C",  -- 76
        58950 => X"38",  -- 56
        58951 => X"42",  -- 66
        58952 => X"2C",  -- 44
        58953 => X"2A",  -- 42
        58954 => X"51",  -- 81
        58955 => X"61",  -- 97
        58956 => X"5C",  -- 92
        58957 => X"52",  -- 82
        58958 => X"7B",  -- 123
        58959 => X"97",  -- 151
        58960 => X"85",  -- 133
        58961 => X"82",  -- 130
        58962 => X"91",  -- 145
        58963 => X"89",  -- 137
        58964 => X"85",  -- 133
        58965 => X"80",  -- 128
        58966 => X"85",  -- 133
        58967 => X"72",  -- 114
        58968 => X"59",  -- 89
        58969 => X"29",  -- 41
        58970 => X"0D",  -- 13
        58971 => X"0F",  -- 15
        58972 => X"0D",  -- 13
        58973 => X"06",  -- 6
        58974 => X"0B",  -- 11
        58975 => X"16",  -- 22
        58976 => X"1A",  -- 26
        58977 => X"49",  -- 73
        58978 => X"83",  -- 131
        58979 => X"7D",  -- 125
        58980 => X"8B",  -- 139
        58981 => X"93",  -- 147
        58982 => X"9F",  -- 159
        58983 => X"99",  -- 153
        58984 => X"A9",  -- 169
        58985 => X"9D",  -- 157
        58986 => X"B5",  -- 181
        58987 => X"97",  -- 151
        58988 => X"81",  -- 129
        58989 => X"99",  -- 153
        58990 => X"81",  -- 129
        58991 => X"64",  -- 100
        58992 => X"5F",  -- 95
        58993 => X"74",  -- 116
        58994 => X"8B",  -- 139
        58995 => X"59",  -- 89
        58996 => X"2C",  -- 44
        58997 => X"43",  -- 67
        58998 => X"72",  -- 114
        58999 => X"A1",  -- 161
        59000 => X"AE",  -- 174
        59001 => X"AE",  -- 174
        59002 => X"B9",  -- 185
        59003 => X"B0",  -- 176
        59004 => X"99",  -- 153
        59005 => X"9C",  -- 156
        59006 => X"A3",  -- 163
        59007 => X"8E",  -- 142
        59008 => X"88",  -- 136
        59009 => X"A7",  -- 167
        59010 => X"83",  -- 131
        59011 => X"A4",  -- 164
        59012 => X"87",  -- 135
        59013 => X"65",  -- 101
        59014 => X"3B",  -- 59
        59015 => X"1A",  -- 26
        59016 => X"1F",  -- 31
        59017 => X"72",  -- 114
        59018 => X"7F",  -- 127
        59019 => X"44",  -- 68
        59020 => X"19",  -- 25
        59021 => X"3B",  -- 59
        59022 => X"8C",  -- 140
        59023 => X"6F",  -- 111
        59024 => X"3F",  -- 63
        59025 => X"64",  -- 100
        59026 => X"38",  -- 56
        59027 => X"29",  -- 41
        59028 => X"5A",  -- 90
        59029 => X"20",  -- 32
        59030 => X"2C",  -- 44
        59031 => X"32",  -- 50
        59032 => X"36",  -- 54
        59033 => X"3A",  -- 58
        59034 => X"37",  -- 55
        59035 => X"35",  -- 53
        59036 => X"46",  -- 70
        59037 => X"66",  -- 102
        59038 => X"7A",  -- 122
        59039 => X"79",  -- 121
        59040 => X"41",  -- 65
        59041 => X"2A",  -- 42
        59042 => X"2C",  -- 44
        59043 => X"3B",  -- 59
        59044 => X"2F",  -- 47
        59045 => X"2A",  -- 42
        59046 => X"30",  -- 48
        59047 => X"1F",  -- 31
        59048 => X"2A",  -- 42
        59049 => X"3C",  -- 60
        59050 => X"45",  -- 69
        59051 => X"62",  -- 98
        59052 => X"40",  -- 64
        59053 => X"2F",  -- 47
        59054 => X"2F",  -- 47
        59055 => X"29",  -- 41
        59056 => X"2C",  -- 44
        59057 => X"31",  -- 49
        59058 => X"35",  -- 53
        59059 => X"3B",  -- 59
        59060 => X"44",  -- 68
        59061 => X"4E",  -- 78
        59062 => X"52",  -- 82
        59063 => X"50",  -- 80
        59064 => X"51",  -- 81
        59065 => X"4A",  -- 74
        59066 => X"47",  -- 71
        59067 => X"47",  -- 71
        59068 => X"42",  -- 66
        59069 => X"42",  -- 66
        59070 => X"58",  -- 88
        59071 => X"73",  -- 115
        59072 => X"76",  -- 118
        59073 => X"67",  -- 103
        59074 => X"5A",  -- 90
        59075 => X"5E",  -- 94
        59076 => X"70",  -- 112
        59077 => X"7B",  -- 123
        59078 => X"75",  -- 117
        59079 => X"67",  -- 103
        59080 => X"5A",  -- 90
        59081 => X"60",  -- 96
        59082 => X"5C",  -- 92
        59083 => X"4F",  -- 79
        59084 => X"45",  -- 69
        59085 => X"44",  -- 68
        59086 => X"41",  -- 65
        59087 => X"3B",  -- 59
        59088 => X"37",  -- 55
        59089 => X"30",  -- 48
        59090 => X"36",  -- 54
        59091 => X"31",  -- 49
        59092 => X"46",  -- 70
        59093 => X"70",  -- 112
        59094 => X"7B",  -- 123
        59095 => X"87",  -- 135
        59096 => X"96",  -- 150
        59097 => X"83",  -- 131
        59098 => X"8E",  -- 142
        59099 => X"96",  -- 150
        59100 => X"8A",  -- 138
        59101 => X"9F",  -- 159
        59102 => X"BD",  -- 189
        59103 => X"B7",  -- 183
        59104 => X"A1",  -- 161
        59105 => X"8B",  -- 139
        59106 => X"71",  -- 113
        59107 => X"4D",  -- 77
        59108 => X"54",  -- 84
        59109 => X"6E",  -- 110
        59110 => X"73",  -- 115
        59111 => X"8C",  -- 140
        59112 => X"9A",  -- 154
        59113 => X"9B",  -- 155
        59114 => X"B3",  -- 179
        59115 => X"AE",  -- 174
        59116 => X"B3",  -- 179
        59117 => X"AE",  -- 174
        59118 => X"A4",  -- 164
        59119 => X"7A",  -- 122
        59120 => X"85",  -- 133
        59121 => X"8D",  -- 141
        59122 => X"8F",  -- 143
        59123 => X"AF",  -- 175
        59124 => X"AB",  -- 171
        59125 => X"C2",  -- 194
        59126 => X"AF",  -- 175
        59127 => X"B6",  -- 182
        59128 => X"AA",  -- 170
        59129 => X"A5",  -- 165
        59130 => X"A9",  -- 169
        59131 => X"B7",  -- 183
        59132 => X"C1",  -- 193
        59133 => X"BC",  -- 188
        59134 => X"B7",  -- 183
        59135 => X"B5",  -- 181
        59136 => X"A2",  -- 162
        59137 => X"B9",  -- 185
        59138 => X"D9",  -- 217
        59139 => X"A8",  -- 168
        59140 => X"82",  -- 130
        59141 => X"AB",  -- 171
        59142 => X"C3",  -- 195
        59143 => X"C1",  -- 193
        59144 => X"BF",  -- 191
        59145 => X"B9",  -- 185
        59146 => X"BF",  -- 191
        59147 => X"C6",  -- 198
        59148 => X"C2",  -- 194
        59149 => X"C2",  -- 194
        59150 => X"C2",  -- 194
        59151 => X"C0",  -- 192
        59152 => X"CB",  -- 203
        59153 => X"C8",  -- 200
        59154 => X"8E",  -- 142
        59155 => X"36",  -- 54
        59156 => X"1F",  -- 31
        59157 => X"23",  -- 35
        59158 => X"43",  -- 67
        59159 => X"36",  -- 54
        59160 => X"3E",  -- 62
        59161 => X"35",  -- 53
        59162 => X"27",  -- 39
        59163 => X"26",  -- 38
        59164 => X"2E",  -- 46
        59165 => X"2C",  -- 44
        59166 => X"2C",  -- 44
        59167 => X"36",  -- 54
        59168 => X"25",  -- 37
        59169 => X"20",  -- 32
        59170 => X"21",  -- 33
        59171 => X"28",  -- 40
        59172 => X"28",  -- 40
        59173 => X"1E",  -- 30
        59174 => X"15",  -- 21
        59175 => X"13",  -- 19
        59176 => X"1E",  -- 30
        59177 => X"18",  -- 24
        59178 => X"17",  -- 23
        59179 => X"1D",  -- 29
        59180 => X"24",  -- 36
        59181 => X"2A",  -- 42
        59182 => X"33",  -- 51
        59183 => X"3C",  -- 60
        59184 => X"39",  -- 57
        59185 => X"3E",  -- 62
        59186 => X"44",  -- 68
        59187 => X"46",  -- 70
        59188 => X"49",  -- 73
        59189 => X"50",  -- 80
        59190 => X"58",  -- 88
        59191 => X"5C",  -- 92
        59192 => X"60",  -- 96
        59193 => X"6A",  -- 106
        59194 => X"6E",  -- 110
        59195 => X"6E",  -- 110
        59196 => X"75",  -- 117
        59197 => X"7A",  -- 122
        59198 => X"83",  -- 131
        59199 => X"91",  -- 145
        59200 => X"25",  -- 37
        59201 => X"27",  -- 39
        59202 => X"29",  -- 41
        59203 => X"2A",  -- 42
        59204 => X"2F",  -- 47
        59205 => X"35",  -- 53
        59206 => X"34",  -- 52
        59207 => X"2F",  -- 47
        59208 => X"29",  -- 41
        59209 => X"2B",  -- 43
        59210 => X"2D",  -- 45
        59211 => X"29",  -- 41
        59212 => X"24",  -- 36
        59213 => X"1F",  -- 31
        59214 => X"21",  -- 33
        59215 => X"25",  -- 37
        59216 => X"27",  -- 39
        59217 => X"24",  -- 36
        59218 => X"1D",  -- 29
        59219 => X"1D",  -- 29
        59220 => X"24",  -- 36
        59221 => X"2D",  -- 45
        59222 => X"2E",  -- 46
        59223 => X"27",  -- 39
        59224 => X"3D",  -- 61
        59225 => X"34",  -- 52
        59226 => X"3E",  -- 62
        59227 => X"38",  -- 56
        59228 => X"31",  -- 49
        59229 => X"36",  -- 54
        59230 => X"4B",  -- 75
        59231 => X"7F",  -- 127
        59232 => X"5B",  -- 91
        59233 => X"26",  -- 38
        59234 => X"25",  -- 37
        59235 => X"34",  -- 52
        59236 => X"9C",  -- 156
        59237 => X"50",  -- 80
        59238 => X"1E",  -- 30
        59239 => X"21",  -- 33
        59240 => X"2D",  -- 45
        59241 => X"13",  -- 19
        59242 => X"58",  -- 88
        59243 => X"9E",  -- 158
        59244 => X"99",  -- 153
        59245 => X"83",  -- 131
        59246 => X"7A",  -- 122
        59247 => X"81",  -- 129
        59248 => X"2B",  -- 43
        59249 => X"34",  -- 52
        59250 => X"8A",  -- 138
        59251 => X"6A",  -- 106
        59252 => X"2E",  -- 46
        59253 => X"1C",  -- 28
        59254 => X"50",  -- 80
        59255 => X"56",  -- 86
        59256 => X"70",  -- 112
        59257 => X"1B",  -- 27
        59258 => X"21",  -- 33
        59259 => X"53",  -- 83
        59260 => X"46",  -- 70
        59261 => X"61",  -- 97
        59262 => X"64",  -- 100
        59263 => X"3B",  -- 59
        59264 => X"66",  -- 102
        59265 => X"7B",  -- 123
        59266 => X"71",  -- 113
        59267 => X"7F",  -- 127
        59268 => X"97",  -- 151
        59269 => X"71",  -- 113
        59270 => X"52",  -- 82
        59271 => X"6C",  -- 108
        59272 => X"58",  -- 88
        59273 => X"42",  -- 66
        59274 => X"45",  -- 69
        59275 => X"3D",  -- 61
        59276 => X"2F",  -- 47
        59277 => X"23",  -- 35
        59278 => X"49",  -- 73
        59279 => X"67",  -- 103
        59280 => X"49",  -- 73
        59281 => X"59",  -- 89
        59282 => X"71",  -- 113
        59283 => X"6F",  -- 111
        59284 => X"76",  -- 118
        59285 => X"6E",  -- 110
        59286 => X"78",  -- 120
        59287 => X"7A",  -- 122
        59288 => X"70",  -- 112
        59289 => X"4B",  -- 75
        59290 => X"25",  -- 37
        59291 => X"16",  -- 22
        59292 => X"0C",  -- 12
        59293 => X"03",  -- 3
        59294 => X"0E",  -- 14
        59295 => X"23",  -- 35
        59296 => X"54",  -- 84
        59297 => X"73",  -- 115
        59298 => X"84",  -- 132
        59299 => X"89",  -- 137
        59300 => X"78",  -- 120
        59301 => X"85",  -- 133
        59302 => X"7C",  -- 124
        59303 => X"7C",  -- 124
        59304 => X"7A",  -- 122
        59305 => X"69",  -- 105
        59306 => X"6D",  -- 109
        59307 => X"4B",  -- 75
        59308 => X"33",  -- 51
        59309 => X"49",  -- 73
        59310 => X"46",  -- 70
        59311 => X"35",  -- 53
        59312 => X"38",  -- 56
        59313 => X"5E",  -- 94
        59314 => X"83",  -- 131
        59315 => X"78",  -- 120
        59316 => X"69",  -- 105
        59317 => X"82",  -- 130
        59318 => X"A4",  -- 164
        59319 => X"B9",  -- 185
        59320 => X"CB",  -- 203
        59321 => X"BB",  -- 187
        59322 => X"AE",  -- 174
        59323 => X"96",  -- 150
        59324 => X"7C",  -- 124
        59325 => X"82",  -- 130
        59326 => X"97",  -- 151
        59327 => X"9B",  -- 155
        59328 => X"9A",  -- 154
        59329 => X"B0",  -- 176
        59330 => X"7F",  -- 127
        59331 => X"7A",  -- 122
        59332 => X"7E",  -- 126
        59333 => X"A9",  -- 169
        59334 => X"CA",  -- 202
        59335 => X"7D",  -- 125
        59336 => X"3F",  -- 63
        59337 => X"0C",  -- 12
        59338 => X"50",  -- 80
        59339 => X"8F",  -- 143
        59340 => X"7B",  -- 123
        59341 => X"26",  -- 38
        59342 => X"1A",  -- 26
        59343 => X"61",  -- 97
        59344 => X"83",  -- 131
        59345 => X"47",  -- 71
        59346 => X"55",  -- 85
        59347 => X"4A",  -- 74
        59348 => X"38",  -- 56
        59349 => X"41",  -- 65
        59350 => X"26",  -- 38
        59351 => X"38",  -- 56
        59352 => X"38",  -- 56
        59353 => X"48",  -- 72
        59354 => X"36",  -- 54
        59355 => X"2A",  -- 42
        59356 => X"37",  -- 55
        59357 => X"34",  -- 52
        59358 => X"43",  -- 67
        59359 => X"79",  -- 121
        59360 => X"8A",  -- 138
        59361 => X"5A",  -- 90
        59362 => X"3E",  -- 62
        59363 => X"32",  -- 50
        59364 => X"37",  -- 55
        59365 => X"3A",  -- 58
        59366 => X"2B",  -- 43
        59367 => X"37",  -- 55
        59368 => X"3C",  -- 60
        59369 => X"3D",  -- 61
        59370 => X"2C",  -- 44
        59371 => X"3F",  -- 63
        59372 => X"36",  -- 54
        59373 => X"35",  -- 53
        59374 => X"32",  -- 50
        59375 => X"28",  -- 40
        59376 => X"2A",  -- 42
        59377 => X"33",  -- 51
        59378 => X"3B",  -- 59
        59379 => X"3B",  -- 59
        59380 => X"3C",  -- 60
        59381 => X"44",  -- 68
        59382 => X"4F",  -- 79
        59383 => X"56",  -- 86
        59384 => X"47",  -- 71
        59385 => X"3F",  -- 63
        59386 => X"3B",  -- 59
        59387 => X"3E",  -- 62
        59388 => X"3E",  -- 62
        59389 => X"40",  -- 64
        59390 => X"54",  -- 84
        59391 => X"6C",  -- 108
        59392 => X"6F",  -- 111
        59393 => X"65",  -- 101
        59394 => X"5A",  -- 90
        59395 => X"5A",  -- 90
        59396 => X"68",  -- 104
        59397 => X"72",  -- 114
        59398 => X"6D",  -- 109
        59399 => X"63",  -- 99
        59400 => X"5B",  -- 91
        59401 => X"61",  -- 97
        59402 => X"60",  -- 96
        59403 => X"53",  -- 83
        59404 => X"4B",  -- 75
        59405 => X"48",  -- 72
        59406 => X"45",  -- 69
        59407 => X"3E",  -- 62
        59408 => X"3B",  -- 59
        59409 => X"33",  -- 51
        59410 => X"38",  -- 56
        59411 => X"37",  -- 55
        59412 => X"50",  -- 80
        59413 => X"79",  -- 121
        59414 => X"86",  -- 134
        59415 => X"90",  -- 144
        59416 => X"8D",  -- 141
        59417 => X"87",  -- 135
        59418 => X"90",  -- 144
        59419 => X"97",  -- 151
        59420 => X"98",  -- 152
        59421 => X"AA",  -- 170
        59422 => X"AF",  -- 175
        59423 => X"97",  -- 151
        59424 => X"84",  -- 132
        59425 => X"69",  -- 105
        59426 => X"5D",  -- 93
        59427 => X"53",  -- 83
        59428 => X"57",  -- 87
        59429 => X"79",  -- 121
        59430 => X"96",  -- 150
        59431 => X"A5",  -- 165
        59432 => X"96",  -- 150
        59433 => X"A7",  -- 167
        59434 => X"BA",  -- 186
        59435 => X"A7",  -- 167
        59436 => X"A4",  -- 164
        59437 => X"A9",  -- 169
        59438 => X"A9",  -- 169
        59439 => X"70",  -- 112
        59440 => X"8C",  -- 140
        59441 => X"8F",  -- 143
        59442 => X"98",  -- 152
        59443 => X"B8",  -- 184
        59444 => X"B6",  -- 182
        59445 => X"BC",  -- 188
        59446 => X"B1",  -- 177
        59447 => X"C7",  -- 199
        59448 => X"C1",  -- 193
        59449 => X"C2",  -- 194
        59450 => X"C0",  -- 192
        59451 => X"BD",  -- 189
        59452 => X"BB",  -- 187
        59453 => X"BE",  -- 190
        59454 => X"BD",  -- 189
        59455 => X"BC",  -- 188
        59456 => X"B5",  -- 181
        59457 => X"BC",  -- 188
        59458 => X"CF",  -- 207
        59459 => X"A7",  -- 167
        59460 => X"88",  -- 136
        59461 => X"A3",  -- 163
        59462 => X"BB",  -- 187
        59463 => X"CC",  -- 204
        59464 => X"CD",  -- 205
        59465 => X"C2",  -- 194
        59466 => X"C2",  -- 194
        59467 => X"C3",  -- 195
        59468 => X"BC",  -- 188
        59469 => X"BD",  -- 189
        59470 => X"C3",  -- 195
        59471 => X"C3",  -- 195
        59472 => X"C0",  -- 192
        59473 => X"C9",  -- 201
        59474 => X"B8",  -- 184
        59475 => X"60",  -- 96
        59476 => X"21",  -- 33
        59477 => X"21",  -- 33
        59478 => X"32",  -- 50
        59479 => X"31",  -- 49
        59480 => X"3B",  -- 59
        59481 => X"33",  -- 51
        59482 => X"28",  -- 40
        59483 => X"26",  -- 38
        59484 => X"2C",  -- 44
        59485 => X"2A",  -- 42
        59486 => X"29",  -- 41
        59487 => X"33",  -- 51
        59488 => X"28",  -- 40
        59489 => X"20",  -- 32
        59490 => X"1D",  -- 29
        59491 => X"24",  -- 36
        59492 => X"29",  -- 41
        59493 => X"21",  -- 33
        59494 => X"17",  -- 23
        59495 => X"13",  -- 19
        59496 => X"19",  -- 25
        59497 => X"15",  -- 21
        59498 => X"16",  -- 22
        59499 => X"1D",  -- 29
        59500 => X"24",  -- 36
        59501 => X"29",  -- 41
        59502 => X"31",  -- 49
        59503 => X"38",  -- 56
        59504 => X"3B",  -- 59
        59505 => X"41",  -- 65
        59506 => X"45",  -- 69
        59507 => X"49",  -- 73
        59508 => X"4E",  -- 78
        59509 => X"58",  -- 88
        59510 => X"60",  -- 96
        59511 => X"63",  -- 99
        59512 => X"69",  -- 105
        59513 => X"72",  -- 114
        59514 => X"73",  -- 115
        59515 => X"72",  -- 114
        59516 => X"77",  -- 119
        59517 => X"7C",  -- 124
        59518 => X"85",  -- 133
        59519 => X"93",  -- 147
        59520 => X"32",  -- 50
        59521 => X"32",  -- 50
        59522 => X"32",  -- 50
        59523 => X"34",  -- 52
        59524 => X"38",  -- 56
        59525 => X"3A",  -- 58
        59526 => X"33",  -- 51
        59527 => X"2A",  -- 42
        59528 => X"22",  -- 34
        59529 => X"27",  -- 39
        59530 => X"2B",  -- 43
        59531 => X"26",  -- 38
        59532 => X"1F",  -- 31
        59533 => X"1A",  -- 26
        59534 => X"1D",  -- 29
        59535 => X"21",  -- 33
        59536 => X"2C",  -- 44
        59537 => X"2D",  -- 45
        59538 => X"26",  -- 38
        59539 => X"1F",  -- 31
        59540 => X"26",  -- 38
        59541 => X"33",  -- 51
        59542 => X"34",  -- 52
        59543 => X"2D",  -- 45
        59544 => X"2A",  -- 42
        59545 => X"40",  -- 64
        59546 => X"43",  -- 67
        59547 => X"3C",  -- 60
        59548 => X"33",  -- 51
        59549 => X"63",  -- 99
        59550 => X"8D",  -- 141
        59551 => X"48",  -- 72
        59552 => X"2B",  -- 43
        59553 => X"26",  -- 38
        59554 => X"2C",  -- 44
        59555 => X"79",  -- 121
        59556 => X"4D",  -- 77
        59557 => X"22",  -- 34
        59558 => X"19",  -- 25
        59559 => X"38",  -- 56
        59560 => X"2A",  -- 42
        59561 => X"64",  -- 100
        59562 => X"AB",  -- 171
        59563 => X"9B",  -- 155
        59564 => X"7F",  -- 127
        59565 => X"89",  -- 137
        59566 => X"5A",  -- 90
        59567 => X"14",  -- 20
        59568 => X"34",  -- 52
        59569 => X"8A",  -- 138
        59570 => X"54",  -- 84
        59571 => X"25",  -- 37
        59572 => X"24",  -- 36
        59573 => X"5E",  -- 94
        59574 => X"68",  -- 104
        59575 => X"5A",  -- 90
        59576 => X"1A",  -- 26
        59577 => X"2C",  -- 44
        59578 => X"62",  -- 98
        59579 => X"33",  -- 51
        59580 => X"70",  -- 112
        59581 => X"74",  -- 116
        59582 => X"57",  -- 87
        59583 => X"47",  -- 71
        59584 => X"4E",  -- 78
        59585 => X"47",  -- 71
        59586 => X"4E",  -- 78
        59587 => X"78",  -- 120
        59588 => X"79",  -- 121
        59589 => X"73",  -- 115
        59590 => X"94",  -- 148
        59591 => X"8E",  -- 142
        59592 => X"87",  -- 135
        59593 => X"70",  -- 112
        59594 => X"67",  -- 103
        59595 => X"56",  -- 86
        59596 => X"58",  -- 88
        59597 => X"58",  -- 88
        59598 => X"6C",  -- 108
        59599 => X"6B",  -- 107
        59600 => X"6A",  -- 106
        59601 => X"68",  -- 104
        59602 => X"67",  -- 103
        59603 => X"60",  -- 96
        59604 => X"74",  -- 116
        59605 => X"71",  -- 113
        59606 => X"7D",  -- 125
        59607 => X"88",  -- 136
        59608 => X"72",  -- 114
        59609 => X"6D",  -- 109
        59610 => X"50",  -- 80
        59611 => X"2E",  -- 46
        59612 => X"18",  -- 24
        59613 => X"0A",  -- 10
        59614 => X"1B",  -- 27
        59615 => X"43",  -- 67
        59616 => X"61",  -- 97
        59617 => X"71",  -- 113
        59618 => X"75",  -- 117
        59619 => X"83",  -- 131
        59620 => X"73",  -- 115
        59621 => X"75",  -- 117
        59622 => X"69",  -- 105
        59623 => X"6B",  -- 107
        59624 => X"72",  -- 114
        59625 => X"69",  -- 105
        59626 => X"75",  -- 117
        59627 => X"7D",  -- 125
        59628 => X"82",  -- 130
        59629 => X"8E",  -- 142
        59630 => X"84",  -- 132
        59631 => X"64",  -- 100
        59632 => X"6A",  -- 106
        59633 => X"87",  -- 135
        59634 => X"A2",  -- 162
        59635 => X"B3",  -- 179
        59636 => X"B2",  -- 178
        59637 => X"B2",  -- 178
        59638 => X"AD",  -- 173
        59639 => X"91",  -- 145
        59640 => X"AC",  -- 172
        59641 => X"8F",  -- 143
        59642 => X"82",  -- 130
        59643 => X"8D",  -- 141
        59644 => X"8C",  -- 140
        59645 => X"72",  -- 114
        59646 => X"57",  -- 87
        59647 => X"4B",  -- 75
        59648 => X"53",  -- 83
        59649 => X"72",  -- 114
        59650 => X"D2",  -- 210
        59651 => X"9C",  -- 156
        59652 => X"68",  -- 104
        59653 => X"88",  -- 136
        59654 => X"8A",  -- 138
        59655 => X"8F",  -- 143
        59656 => X"99",  -- 153
        59657 => X"8B",  -- 139
        59658 => X"3C",  -- 60
        59659 => X"4B",  -- 75
        59660 => X"43",  -- 67
        59661 => X"7F",  -- 127
        59662 => X"68",  -- 104
        59663 => X"24",  -- 36
        59664 => X"37",  -- 55
        59665 => X"A2",  -- 162
        59666 => X"61",  -- 97
        59667 => X"3C",  -- 60
        59668 => X"6C",  -- 108
        59669 => X"59",  -- 89
        59670 => X"3A",  -- 58
        59671 => X"35",  -- 53
        59672 => X"38",  -- 56
        59673 => X"2F",  -- 47
        59674 => X"3B",  -- 59
        59675 => X"47",  -- 71
        59676 => X"37",  -- 55
        59677 => X"29",  -- 41
        59678 => X"31",  -- 49
        59679 => X"3E",  -- 62
        59680 => X"56",  -- 86
        59681 => X"8C",  -- 140
        59682 => X"5D",  -- 93
        59683 => X"37",  -- 55
        59684 => X"40",  -- 64
        59685 => X"32",  -- 50
        59686 => X"2D",  -- 45
        59687 => X"2C",  -- 44
        59688 => X"32",  -- 50
        59689 => X"3E",  -- 62
        59690 => X"32",  -- 50
        59691 => X"35",  -- 53
        59692 => X"31",  -- 49
        59693 => X"2F",  -- 47
        59694 => X"2B",  -- 43
        59695 => X"2A",  -- 42
        59696 => X"2A",  -- 42
        59697 => X"30",  -- 48
        59698 => X"33",  -- 51
        59699 => X"31",  -- 49
        59700 => X"33",  -- 51
        59701 => X"3D",  -- 61
        59702 => X"49",  -- 73
        59703 => X"50",  -- 80
        59704 => X"45",  -- 69
        59705 => X"3B",  -- 59
        59706 => X"34",  -- 52
        59707 => X"36",  -- 54
        59708 => X"37",  -- 55
        59709 => X"38",  -- 56
        59710 => X"46",  -- 70
        59711 => X"58",  -- 88
        59712 => X"65",  -- 101
        59713 => X"62",  -- 98
        59714 => X"5C",  -- 92
        59715 => X"59",  -- 89
        59716 => X"5E",  -- 94
        59717 => X"64",  -- 100
        59718 => X"63",  -- 99
        59719 => X"5C",  -- 92
        59720 => X"59",  -- 89
        59721 => X"5E",  -- 94
        59722 => X"5C",  -- 92
        59723 => X"51",  -- 81
        59724 => X"49",  -- 73
        59725 => X"45",  -- 69
        59726 => X"41",  -- 65
        59727 => X"3A",  -- 58
        59728 => X"3A",  -- 58
        59729 => X"31",  -- 49
        59730 => X"34",  -- 52
        59731 => X"3B",  -- 59
        59732 => X"59",  -- 89
        59733 => X"80",  -- 128
        59734 => X"8C",  -- 140
        59735 => X"94",  -- 148
        59736 => X"92",  -- 146
        59737 => X"95",  -- 149
        59738 => X"9A",  -- 154
        59739 => X"9D",  -- 157
        59740 => X"AB",  -- 171
        59741 => X"B3",  -- 179
        59742 => X"9E",  -- 158
        59743 => X"7B",  -- 123
        59744 => X"67",  -- 103
        59745 => X"50",  -- 80
        59746 => X"55",  -- 85
        59747 => X"69",  -- 105
        59748 => X"65",  -- 101
        59749 => X"7A",  -- 122
        59750 => X"A3",  -- 163
        59751 => X"A3",  -- 163
        59752 => X"A1",  -- 161
        59753 => X"B3",  -- 179
        59754 => X"B9",  -- 185
        59755 => X"AC",  -- 172
        59756 => X"A2",  -- 162
        59757 => X"A4",  -- 164
        59758 => X"AA",  -- 170
        59759 => X"6D",  -- 109
        59760 => X"90",  -- 144
        59761 => X"92",  -- 146
        59762 => X"97",  -- 151
        59763 => X"B1",  -- 177
        59764 => X"BE",  -- 190
        59765 => X"BE",  -- 190
        59766 => X"BA",  -- 186
        59767 => X"C9",  -- 201
        59768 => X"C8",  -- 200
        59769 => X"CF",  -- 207
        59770 => X"CF",  -- 207
        59771 => X"C1",  -- 193
        59772 => X"BA",  -- 186
        59773 => X"C0",  -- 192
        59774 => X"C3",  -- 195
        59775 => X"C1",  -- 193
        59776 => X"C6",  -- 198
        59777 => X"C1",  -- 193
        59778 => X"C6",  -- 198
        59779 => X"A2",  -- 162
        59780 => X"8F",  -- 143
        59781 => X"A2",  -- 162
        59782 => X"B2",  -- 178
        59783 => X"D1",  -- 209
        59784 => X"D4",  -- 212
        59785 => X"C8",  -- 200
        59786 => X"C5",  -- 197
        59787 => X"C3",  -- 195
        59788 => X"BC",  -- 188
        59789 => X"BE",  -- 190
        59790 => X"C6",  -- 198
        59791 => X"C8",  -- 200
        59792 => X"BF",  -- 191
        59793 => X"C9",  -- 201
        59794 => X"D9",  -- 217
        59795 => X"90",  -- 144
        59796 => X"2C",  -- 44
        59797 => X"25",  -- 37
        59798 => X"27",  -- 39
        59799 => X"2D",  -- 45
        59800 => X"35",  -- 53
        59801 => X"30",  -- 48
        59802 => X"29",  -- 41
        59803 => X"2A",  -- 42
        59804 => X"2D",  -- 45
        59805 => X"27",  -- 39
        59806 => X"25",  -- 37
        59807 => X"31",  -- 49
        59808 => X"2D",  -- 45
        59809 => X"1F",  -- 31
        59810 => X"18",  -- 24
        59811 => X"20",  -- 32
        59812 => X"28",  -- 40
        59813 => X"25",  -- 37
        59814 => X"1A",  -- 26
        59815 => X"14",  -- 20
        59816 => X"17",  -- 23
        59817 => X"16",  -- 22
        59818 => X"18",  -- 24
        59819 => X"1E",  -- 30
        59820 => X"25",  -- 37
        59821 => X"2A",  -- 42
        59822 => X"31",  -- 49
        59823 => X"36",  -- 54
        59824 => X"3D",  -- 61
        59825 => X"44",  -- 68
        59826 => X"48",  -- 72
        59827 => X"4D",  -- 77
        59828 => X"58",  -- 88
        59829 => X"64",  -- 100
        59830 => X"6C",  -- 108
        59831 => X"6D",  -- 109
        59832 => X"73",  -- 115
        59833 => X"7B",  -- 123
        59834 => X"79",  -- 121
        59835 => X"77",  -- 119
        59836 => X"7C",  -- 124
        59837 => X"80",  -- 128
        59838 => X"88",  -- 136
        59839 => X"95",  -- 149
        59840 => X"53",  -- 83
        59841 => X"53",  -- 83
        59842 => X"53",  -- 83
        59843 => X"4F",  -- 79
        59844 => X"4E",  -- 78
        59845 => X"4D",  -- 77
        59846 => X"46",  -- 70
        59847 => X"3E",  -- 62
        59848 => X"3C",  -- 60
        59849 => X"3E",  -- 62
        59850 => X"3F",  -- 63
        59851 => X"3C",  -- 60
        59852 => X"35",  -- 53
        59853 => X"2E",  -- 46
        59854 => X"2C",  -- 44
        59855 => X"2C",  -- 44
        59856 => X"36",  -- 54
        59857 => X"36",  -- 54
        59858 => X"2E",  -- 46
        59859 => X"28",  -- 40
        59860 => X"30",  -- 48
        59861 => X"3E",  -- 62
        59862 => X"3D",  -- 61
        59863 => X"30",  -- 48
        59864 => X"3D",  -- 61
        59865 => X"3E",  -- 62
        59866 => X"42",  -- 66
        59867 => X"3B",  -- 59
        59868 => X"6B",  -- 107
        59869 => X"7F",  -- 127
        59870 => X"41",  -- 65
        59871 => X"35",  -- 53
        59872 => X"2A",  -- 42
        59873 => X"2F",  -- 47
        59874 => X"80",  -- 128
        59875 => X"73",  -- 115
        59876 => X"26",  -- 38
        59877 => X"24",  -- 36
        59878 => X"1D",  -- 29
        59879 => X"49",  -- 73
        59880 => X"8E",  -- 142
        59881 => X"AD",  -- 173
        59882 => X"71",  -- 113
        59883 => X"74",  -- 116
        59884 => X"64",  -- 100
        59885 => X"21",  -- 33
        59886 => X"2E",  -- 46
        59887 => X"2C",  -- 44
        59888 => X"6B",  -- 107
        59889 => X"4C",  -- 76
        59890 => X"27",  -- 39
        59891 => X"12",  -- 18
        59892 => X"71",  -- 113
        59893 => X"97",  -- 151
        59894 => X"48",  -- 72
        59895 => X"18",  -- 24
        59896 => X"32",  -- 50
        59897 => X"58",  -- 88
        59898 => X"34",  -- 52
        59899 => X"8A",  -- 138
        59900 => X"7E",  -- 126
        59901 => X"3C",  -- 60
        59902 => X"3F",  -- 63
        59903 => X"4D",  -- 77
        59904 => X"49",  -- 73
        59905 => X"58",  -- 88
        59906 => X"3E",  -- 62
        59907 => X"31",  -- 49
        59908 => X"41",  -- 65
        59909 => X"53",  -- 83
        59910 => X"6C",  -- 108
        59911 => X"76",  -- 118
        59912 => X"67",  -- 103
        59913 => X"7A",  -- 122
        59914 => X"8F",  -- 143
        59915 => X"84",  -- 132
        59916 => X"8E",  -- 142
        59917 => X"93",  -- 147
        59918 => X"96",  -- 150
        59919 => X"80",  -- 128
        59920 => X"83",  -- 131
        59921 => X"76",  -- 118
        59922 => X"81",  -- 129
        59923 => X"84",  -- 132
        59924 => X"85",  -- 133
        59925 => X"74",  -- 116
        59926 => X"74",  -- 116
        59927 => X"6A",  -- 106
        59928 => X"5F",  -- 95
        59929 => X"77",  -- 119
        59930 => X"69",  -- 105
        59931 => X"42",  -- 66
        59932 => X"24",  -- 36
        59933 => X"14",  -- 20
        59934 => X"28",  -- 40
        59935 => X"5B",  -- 91
        59936 => X"68",  -- 104
        59937 => X"6B",  -- 107
        59938 => X"7A",  -- 122
        59939 => X"7E",  -- 126
        59940 => X"86",  -- 134
        59941 => X"71",  -- 113
        59942 => X"81",  -- 129
        59943 => X"87",  -- 135
        59944 => X"8B",  -- 139
        59945 => X"86",  -- 134
        59946 => X"87",  -- 135
        59947 => X"98",  -- 152
        59948 => X"9D",  -- 157
        59949 => X"9F",  -- 159
        59950 => X"A3",  -- 163
        59951 => X"92",  -- 146
        59952 => X"8E",  -- 142
        59953 => X"9E",  -- 158
        59954 => X"A3",  -- 163
        59955 => X"B1",  -- 177
        59956 => X"A5",  -- 165
        59957 => X"89",  -- 137
        59958 => X"80",  -- 128
        59959 => X"61",  -- 97
        59960 => X"5E",  -- 94
        59961 => X"66",  -- 102
        59962 => X"70",  -- 112
        59963 => X"8A",  -- 138
        59964 => X"A7",  -- 167
        59965 => X"A3",  -- 163
        59966 => X"7E",  -- 126
        59967 => X"5D",  -- 93
        59968 => X"55",  -- 85
        59969 => X"3E",  -- 62
        59970 => X"4D",  -- 77
        59971 => X"87",  -- 135
        59972 => X"BC",  -- 188
        59973 => X"93",  -- 147
        59974 => X"78",  -- 120
        59975 => X"A8",  -- 168
        59976 => X"79",  -- 121
        59977 => X"3E",  -- 62
        59978 => X"86",  -- 134
        59979 => X"8C",  -- 140
        59980 => X"58",  -- 88
        59981 => X"48",  -- 72
        59982 => X"65",  -- 101
        59983 => X"75",  -- 117
        59984 => X"26",  -- 38
        59985 => X"1C",  -- 28
        59986 => X"85",  -- 133
        59987 => X"68",  -- 104
        59988 => X"3A",  -- 58
        59989 => X"62",  -- 98
        59990 => X"7E",  -- 126
        59991 => X"20",  -- 32
        59992 => X"3D",  -- 61
        59993 => X"27",  -- 39
        59994 => X"37",  -- 55
        59995 => X"43",  -- 67
        59996 => X"2C",  -- 44
        59997 => X"32",  -- 50
        59998 => X"3F",  -- 63
        59999 => X"28",  -- 40
        60000 => X"33",  -- 51
        60001 => X"45",  -- 69
        60002 => X"82",  -- 130
        60003 => X"6F",  -- 111
        60004 => X"42",  -- 66
        60005 => X"3D",  -- 61
        60006 => X"28",  -- 40
        60007 => X"1E",  -- 30
        60008 => X"24",  -- 36
        60009 => X"3E",  -- 62
        60010 => X"3D",  -- 61
        60011 => X"37",  -- 55
        60012 => X"33",  -- 51
        60013 => X"2D",  -- 45
        60014 => X"29",  -- 41
        60015 => X"30",  -- 48
        60016 => X"34",  -- 52
        60017 => X"30",  -- 48
        60018 => X"29",  -- 41
        60019 => X"29",  -- 41
        60020 => X"33",  -- 51
        60021 => X"3F",  -- 63
        60022 => X"44",  -- 68
        60023 => X"43",  -- 67
        60024 => X"45",  -- 69
        60025 => X"3D",  -- 61
        60026 => X"38",  -- 56
        60027 => X"36",  -- 54
        60028 => X"33",  -- 51
        60029 => X"32",  -- 50
        60030 => X"3C",  -- 60
        60031 => X"4B",  -- 75
        60032 => X"61",  -- 97
        60033 => X"65",  -- 101
        60034 => X"62",  -- 98
        60035 => X"5B",  -- 91
        60036 => X"58",  -- 88
        60037 => X"5C",  -- 92
        60038 => X"5C",  -- 92
        60039 => X"59",  -- 89
        60040 => X"58",  -- 88
        60041 => X"5B",  -- 91
        60042 => X"55",  -- 85
        60043 => X"4A",  -- 74
        60044 => X"41",  -- 65
        60045 => X"3C",  -- 60
        60046 => X"37",  -- 55
        60047 => X"33",  -- 51
        60048 => X"36",  -- 54
        60049 => X"2D",  -- 45
        60050 => X"30",  -- 48
        60051 => X"40",  -- 64
        60052 => X"63",  -- 99
        60053 => X"84",  -- 132
        60054 => X"93",  -- 147
        60055 => X"96",  -- 150
        60056 => X"9E",  -- 158
        60057 => X"A4",  -- 164
        60058 => X"9B",  -- 155
        60059 => X"9D",  -- 157
        60060 => X"B1",  -- 177
        60061 => X"B1",  -- 177
        60062 => X"90",  -- 144
        60063 => X"76",  -- 118
        60064 => X"56",  -- 86
        60065 => X"57",  -- 87
        60066 => X"64",  -- 100
        60067 => X"89",  -- 137
        60068 => X"85",  -- 133
        60069 => X"80",  -- 128
        60070 => X"9E",  -- 158
        60071 => X"9C",  -- 156
        60072 => X"B0",  -- 176
        60073 => X"B0",  -- 176
        60074 => X"AC",  -- 172
        60075 => X"B6",  -- 182
        60076 => X"AD",  -- 173
        60077 => X"9F",  -- 159
        60078 => X"9C",  -- 156
        60079 => X"68",  -- 104
        60080 => X"90",  -- 144
        60081 => X"92",  -- 146
        60082 => X"8A",  -- 138
        60083 => X"97",  -- 151
        60084 => X"B7",  -- 183
        60085 => X"BC",  -- 188
        60086 => X"BB",  -- 187
        60087 => X"B6",  -- 182
        60088 => X"BB",  -- 187
        60089 => X"C7",  -- 199
        60090 => X"CF",  -- 207
        60091 => X"CC",  -- 204
        60092 => X"C9",  -- 201
        60093 => X"CA",  -- 202
        60094 => X"C8",  -- 200
        60095 => X"C5",  -- 197
        60096 => X"CC",  -- 204
        60097 => X"C9",  -- 201
        60098 => X"C3",  -- 195
        60099 => X"99",  -- 153
        60100 => X"92",  -- 146
        60101 => X"AD",  -- 173
        60102 => X"B3",  -- 179
        60103 => X"C8",  -- 200
        60104 => X"D0",  -- 208
        60105 => X"C7",  -- 199
        60106 => X"C5",  -- 197
        60107 => X"C7",  -- 199
        60108 => X"C2",  -- 194
        60109 => X"C3",  -- 195
        60110 => X"C9",  -- 201
        60111 => X"CA",  -- 202
        60112 => X"CB",  -- 203
        60113 => X"C9",  -- 201
        60114 => X"D7",  -- 215
        60115 => X"B4",  -- 180
        60116 => X"45",  -- 69
        60117 => X"28",  -- 40
        60118 => X"2B",  -- 43
        60119 => X"2F",  -- 47
        60120 => X"31",  -- 49
        60121 => X"30",  -- 48
        60122 => X"2C",  -- 44
        60123 => X"2B",  -- 43
        60124 => X"2D",  -- 45
        60125 => X"25",  -- 37
        60126 => X"23",  -- 35
        60127 => X"2F",  -- 47
        60128 => X"2F",  -- 47
        60129 => X"21",  -- 33
        60130 => X"19",  -- 25
        60131 => X"20",  -- 32
        60132 => X"27",  -- 39
        60133 => X"24",  -- 36
        60134 => X"1D",  -- 29
        60135 => X"19",  -- 25
        60136 => X"1A",  -- 26
        60137 => X"1A",  -- 26
        60138 => X"1C",  -- 28
        60139 => X"21",  -- 33
        60140 => X"26",  -- 38
        60141 => X"2D",  -- 45
        60142 => X"35",  -- 53
        60143 => X"3B",  -- 59
        60144 => X"3E",  -- 62
        60145 => X"47",  -- 71
        60146 => X"4E",  -- 78
        60147 => X"55",  -- 85
        60148 => X"61",  -- 97
        60149 => X"6F",  -- 111
        60150 => X"74",  -- 116
        60151 => X"72",  -- 114
        60152 => X"79",  -- 121
        60153 => X"80",  -- 128
        60154 => X"7E",  -- 126
        60155 => X"7C",  -- 124
        60156 => X"81",  -- 129
        60157 => X"83",  -- 131
        60158 => X"88",  -- 136
        60159 => X"94",  -- 148
        60160 => X"70",  -- 112
        60161 => X"75",  -- 117
        60162 => X"75",  -- 117
        60163 => X"71",  -- 113
        60164 => X"6C",  -- 108
        60165 => X"6C",  -- 108
        60166 => X"6B",  -- 107
        60167 => X"6A",  -- 106
        60168 => X"6A",  -- 106
        60169 => X"68",  -- 104
        60170 => X"68",  -- 104
        60171 => X"67",  -- 103
        60172 => X"65",  -- 101
        60173 => X"5F",  -- 95
        60174 => X"59",  -- 89
        60175 => X"56",  -- 86
        60176 => X"5D",  -- 93
        60177 => X"5B",  -- 91
        60178 => X"52",  -- 82
        60179 => X"4C",  -- 76
        60180 => X"56",  -- 86
        60181 => X"5F",  -- 95
        60182 => X"58",  -- 88
        60183 => X"49",  -- 73
        60184 => X"53",  -- 83
        60185 => X"5C",  -- 92
        60186 => X"51",  -- 81
        60187 => X"78",  -- 120
        60188 => X"7D",  -- 125
        60189 => X"4E",  -- 78
        60190 => X"4B",  -- 75
        60191 => X"48",  -- 72
        60192 => X"3B",  -- 59
        60193 => X"79",  -- 121
        60194 => X"7A",  -- 122
        60195 => X"2D",  -- 45
        60196 => X"3D",  -- 61
        60197 => X"42",  -- 66
        60198 => X"75",  -- 117
        60199 => X"7F",  -- 127
        60200 => X"9A",  -- 154
        60201 => X"7B",  -- 123
        60202 => X"7A",  -- 122
        60203 => X"42",  -- 66
        60204 => X"36",  -- 54
        60205 => X"37",  -- 55
        60206 => X"17",  -- 23
        60207 => X"5F",  -- 95
        60208 => X"49",  -- 73
        60209 => X"23",  -- 35
        60210 => X"18",  -- 24
        60211 => X"6F",  -- 111
        60212 => X"9B",  -- 155
        60213 => X"41",  -- 65
        60214 => X"24",  -- 36
        60215 => X"2E",  -- 46
        60216 => X"5E",  -- 94
        60217 => X"4A",  -- 74
        60218 => X"5F",  -- 95
        60219 => X"8B",  -- 139
        60220 => X"3F",  -- 63
        60221 => X"2C",  -- 44
        60222 => X"37",  -- 55
        60223 => X"48",  -- 72
        60224 => X"68",  -- 104
        60225 => X"64",  -- 100
        60226 => X"51",  -- 81
        60227 => X"2C",  -- 44
        60228 => X"31",  -- 49
        60229 => X"47",  -- 71
        60230 => X"3A",  -- 58
        60231 => X"33",  -- 51
        60232 => X"36",  -- 54
        60233 => X"5A",  -- 90
        60234 => X"81",  -- 129
        60235 => X"7D",  -- 125
        60236 => X"79",  -- 121
        60237 => X"66",  -- 102
        60238 => X"6A",  -- 106
        60239 => X"6A",  -- 106
        60240 => X"7A",  -- 122
        60241 => X"63",  -- 99
        60242 => X"79",  -- 121
        60243 => X"72",  -- 114
        60244 => X"58",  -- 88
        60245 => X"52",  -- 82
        60246 => X"74",  -- 116
        60247 => X"72",  -- 114
        60248 => X"5D",  -- 93
        60249 => X"6D",  -- 109
        60250 => X"58",  -- 88
        60251 => X"30",  -- 48
        60252 => X"1A",  -- 26
        60253 => X"0F",  -- 15
        60254 => X"20",  -- 32
        60255 => X"49",  -- 73
        60256 => X"61",  -- 97
        60257 => X"67",  -- 103
        60258 => X"72",  -- 114
        60259 => X"73",  -- 115
        60260 => X"75",  -- 117
        60261 => X"5B",  -- 91
        60262 => X"7A",  -- 122
        60263 => X"88",  -- 136
        60264 => X"76",  -- 118
        60265 => X"84",  -- 132
        60266 => X"8C",  -- 140
        60267 => X"8A",  -- 138
        60268 => X"71",  -- 113
        60269 => X"63",  -- 99
        60270 => X"7E",  -- 126
        60271 => X"92",  -- 146
        60272 => X"58",  -- 88
        60273 => X"68",  -- 104
        60274 => X"73",  -- 115
        60275 => X"85",  -- 133
        60276 => X"75",  -- 117
        60277 => X"5D",  -- 93
        60278 => X"6C",  -- 108
        60279 => X"6C",  -- 108
        60280 => X"6A",  -- 106
        60281 => X"99",  -- 153
        60282 => X"97",  -- 151
        60283 => X"64",  -- 100
        60284 => X"58",  -- 88
        60285 => X"78",  -- 120
        60286 => X"85",  -- 133
        60287 => X"74",  -- 116
        60288 => X"73",  -- 115
        60289 => X"5E",  -- 94
        60290 => X"63",  -- 99
        60291 => X"6F",  -- 111
        60292 => X"47",  -- 71
        60293 => X"6D",  -- 109
        60294 => X"A8",  -- 168
        60295 => X"89",  -- 137
        60296 => X"A4",  -- 164
        60297 => X"6F",  -- 111
        60298 => X"2F",  -- 47
        60299 => X"3E",  -- 62
        60300 => X"86",  -- 134
        60301 => X"91",  -- 145
        60302 => X"36",  -- 54
        60303 => X"51",  -- 81
        60304 => X"90",  -- 144
        60305 => X"57",  -- 87
        60306 => X"21",  -- 33
        60307 => X"70",  -- 112
        60308 => X"82",  -- 130
        60309 => X"2F",  -- 47
        60310 => X"7F",  -- 127
        60311 => X"62",  -- 98
        60312 => X"32",  -- 50
        60313 => X"37",  -- 55
        60314 => X"34",  -- 52
        60315 => X"32",  -- 50
        60316 => X"38",  -- 56
        60317 => X"33",  -- 51
        60318 => X"2F",  -- 47
        60319 => X"36",  -- 54
        60320 => X"39",  -- 57
        60321 => X"36",  -- 54
        60322 => X"37",  -- 55
        60323 => X"6F",  -- 111
        60324 => X"6D",  -- 109
        60325 => X"2F",  -- 47
        60326 => X"21",  -- 33
        60327 => X"15",  -- 21
        60328 => X"23",  -- 35
        60329 => X"33",  -- 51
        60330 => X"37",  -- 55
        60331 => X"2C",  -- 44
        60332 => X"32",  -- 50
        60333 => X"32",  -- 50
        60334 => X"2E",  -- 46
        60335 => X"36",  -- 54
        60336 => X"3A",  -- 58
        60337 => X"38",  -- 56
        60338 => X"32",  -- 50
        60339 => X"2F",  -- 47
        60340 => X"35",  -- 53
        60341 => X"3D",  -- 61
        60342 => X"40",  -- 64
        60343 => X"3D",  -- 61
        60344 => X"3D",  -- 61
        60345 => X"3D",  -- 61
        60346 => X"3C",  -- 60
        60347 => X"3D",  -- 61
        60348 => X"38",  -- 56
        60349 => X"35",  -- 53
        60350 => X"3E",  -- 62
        60351 => X"4B",  -- 75
        60352 => X"60",  -- 96
        60353 => X"6B",  -- 107
        60354 => X"6D",  -- 109
        60355 => X"64",  -- 100
        60356 => X"5D",  -- 93
        60357 => X"5C",  -- 92
        60358 => X"5B",  -- 91
        60359 => X"55",  -- 85
        60360 => X"59",  -- 89
        60361 => X"57",  -- 87
        60362 => X"4C",  -- 76
        60363 => X"40",  -- 64
        60364 => X"36",  -- 54
        60365 => X"32",  -- 50
        60366 => X"31",  -- 49
        60367 => X"2F",  -- 47
        60368 => X"31",  -- 49
        60369 => X"2D",  -- 45
        60370 => X"2F",  -- 47
        60371 => X"4A",  -- 74
        60372 => X"6F",  -- 111
        60373 => X"8A",  -- 138
        60374 => X"98",  -- 152
        60375 => X"99",  -- 153
        60376 => X"9F",  -- 159
        60377 => X"A0",  -- 160
        60378 => X"96",  -- 150
        60379 => X"9C",  -- 156
        60380 => X"AE",  -- 174
        60381 => X"A4",  -- 164
        60382 => X"87",  -- 135
        60383 => X"81",  -- 129
        60384 => X"62",  -- 98
        60385 => X"72",  -- 114
        60386 => X"77",  -- 119
        60387 => X"94",  -- 148
        60388 => X"9A",  -- 154
        60389 => X"8A",  -- 138
        60390 => X"9D",  -- 157
        60391 => X"A9",  -- 169
        60392 => X"BA",  -- 186
        60393 => X"B2",  -- 178
        60394 => X"A5",  -- 165
        60395 => X"B7",  -- 183
        60396 => X"B6",  -- 182
        60397 => X"A0",  -- 160
        60398 => X"7F",  -- 127
        60399 => X"4E",  -- 78
        60400 => X"93",  -- 147
        60401 => X"93",  -- 147
        60402 => X"7E",  -- 126
        60403 => X"90",  -- 144
        60404 => X"B0",  -- 176
        60405 => X"AB",  -- 171
        60406 => X"AB",  -- 171
        60407 => X"B0",  -- 176
        60408 => X"BB",  -- 187
        60409 => X"BF",  -- 191
        60410 => X"CA",  -- 202
        60411 => X"D7",  -- 215
        60412 => X"DA",  -- 218
        60413 => X"D2",  -- 210
        60414 => X"CD",  -- 205
        60415 => X"CE",  -- 206
        60416 => X"CF",  -- 207
        60417 => X"D6",  -- 214
        60418 => X"C9",  -- 201
        60419 => X"8D",  -- 141
        60420 => X"89",  -- 137
        60421 => X"BA",  -- 186
        60422 => X"BF",  -- 191
        60423 => X"C1",  -- 193
        60424 => X"CE",  -- 206
        60425 => X"C4",  -- 196
        60426 => X"C4",  -- 196
        60427 => X"C6",  -- 198
        60428 => X"C1",  -- 193
        60429 => X"C3",  -- 195
        60430 => X"CC",  -- 204
        60431 => X"CD",  -- 205
        60432 => X"D1",  -- 209
        60433 => X"CE",  -- 206
        60434 => X"CA",  -- 202
        60435 => X"D1",  -- 209
        60436 => X"6C",  -- 108
        60437 => X"26",  -- 38
        60438 => X"2F",  -- 47
        60439 => X"31",  -- 49
        60440 => X"31",  -- 49
        60441 => X"31",  -- 49
        60442 => X"2D",  -- 45
        60443 => X"2D",  -- 45
        60444 => X"2F",  -- 47
        60445 => X"26",  -- 38
        60446 => X"24",  -- 36
        60447 => X"2E",  -- 46
        60448 => X"2C",  -- 44
        60449 => X"22",  -- 34
        60450 => X"1E",  -- 30
        60451 => X"23",  -- 35
        60452 => X"25",  -- 37
        60453 => X"20",  -- 32
        60454 => X"1D",  -- 29
        60455 => X"1F",  -- 31
        60456 => X"1E",  -- 30
        60457 => X"1F",  -- 31
        60458 => X"20",  -- 32
        60459 => X"21",  -- 33
        60460 => X"26",  -- 38
        60461 => X"2F",  -- 47
        60462 => X"39",  -- 57
        60463 => X"41",  -- 65
        60464 => X"3F",  -- 63
        60465 => X"4C",  -- 76
        60466 => X"57",  -- 87
        60467 => X"5E",  -- 94
        60468 => X"67",  -- 103
        60469 => X"74",  -- 116
        60470 => X"78",  -- 120
        60471 => X"74",  -- 116
        60472 => X"79",  -- 121
        60473 => X"81",  -- 129
        60474 => X"80",  -- 128
        60475 => X"7F",  -- 127
        60476 => X"84",  -- 132
        60477 => X"84",  -- 132
        60478 => X"85",  -- 133
        60479 => X"8E",  -- 142
        60480 => X"6E",  -- 110
        60481 => X"75",  -- 117
        60482 => X"78",  -- 120
        60483 => X"74",  -- 116
        60484 => X"71",  -- 113
        60485 => X"76",  -- 118
        60486 => X"7C",  -- 124
        60487 => X"7F",  -- 127
        60488 => X"78",  -- 120
        60489 => X"77",  -- 119
        60490 => X"76",  -- 118
        60491 => X"79",  -- 121
        60492 => X"7C",  -- 124
        60493 => X"7B",  -- 123
        60494 => X"77",  -- 119
        60495 => X"72",  -- 114
        60496 => X"74",  -- 116
        60497 => X"6E",  -- 110
        60498 => X"68",  -- 104
        60499 => X"68",  -- 104
        60500 => X"6E",  -- 110
        60501 => X"70",  -- 112
        60502 => X"66",  -- 102
        60503 => X"58",  -- 88
        60504 => X"51",  -- 81
        60505 => X"68",  -- 104
        60506 => X"91",  -- 145
        60507 => X"76",  -- 118
        60508 => X"5C",  -- 92
        60509 => X"66",  -- 102
        60510 => X"5D",  -- 93
        60511 => X"62",  -- 98
        60512 => X"94",  -- 148
        60513 => X"7D",  -- 125
        60514 => X"6B",  -- 107
        60515 => X"64",  -- 100
        60516 => X"74",  -- 116
        60517 => X"9E",  -- 158
        60518 => X"67",  -- 103
        60519 => X"61",  -- 97
        60520 => X"8F",  -- 143
        60521 => X"5C",  -- 92
        60522 => X"33",  -- 51
        60523 => X"35",  -- 53
        60524 => X"26",  -- 38
        60525 => X"28",  -- 40
        60526 => X"5B",  -- 91
        60527 => X"69",  -- 105
        60528 => X"32",  -- 50
        60529 => X"23",  -- 35
        60530 => X"6D",  -- 109
        60531 => X"92",  -- 146
        60532 => X"2E",  -- 46
        60533 => X"28",  -- 40
        60534 => X"38",  -- 56
        60535 => X"5A",  -- 90
        60536 => X"49",  -- 73
        60537 => X"41",  -- 65
        60538 => X"99",  -- 153
        60539 => X"3E",  -- 62
        60540 => X"2B",  -- 43
        60541 => X"3A",  -- 58
        60542 => X"4B",  -- 75
        60543 => X"6F",  -- 111
        60544 => X"6F",  -- 111
        60545 => X"3A",  -- 58
        60546 => X"4A",  -- 74
        60547 => X"50",  -- 80
        60548 => X"4B",  -- 75
        60549 => X"67",  -- 103
        60550 => X"5F",  -- 95
        60551 => X"48",  -- 72
        60552 => X"63",  -- 99
        60553 => X"5C",  -- 92
        60554 => X"67",  -- 103
        60555 => X"6E",  -- 110
        60556 => X"70",  -- 112
        60557 => X"4A",  -- 74
        60558 => X"4B",  -- 75
        60559 => X"63",  -- 99
        60560 => X"57",  -- 87
        60561 => X"4A",  -- 74
        60562 => X"6F",  -- 111
        60563 => X"79",  -- 121
        60564 => X"66",  -- 102
        60565 => X"60",  -- 96
        60566 => X"75",  -- 117
        60567 => X"61",  -- 97
        60568 => X"65",  -- 101
        60569 => X"57",  -- 87
        60570 => X"2E",  -- 46
        60571 => X"0A",  -- 10
        60572 => X"03",  -- 3
        60573 => X"05",  -- 5
        60574 => X"0C",  -- 12
        60575 => X"1F",  -- 31
        60576 => X"46",  -- 70
        60577 => X"68",  -- 104
        60578 => X"6C",  -- 108
        60579 => X"8B",  -- 139
        60580 => X"77",  -- 119
        60581 => X"6F",  -- 111
        60582 => X"7C",  -- 124
        60583 => X"86",  -- 134
        60584 => X"54",  -- 84
        60585 => X"69",  -- 105
        60586 => X"81",  -- 129
        60587 => X"7E",  -- 126
        60588 => X"63",  -- 99
        60589 => X"50",  -- 80
        60590 => X"5C",  -- 92
        60591 => X"78",  -- 120
        60592 => X"56",  -- 86
        60593 => X"5D",  -- 93
        60594 => X"6F",  -- 111
        60595 => X"8E",  -- 142
        60596 => X"94",  -- 148
        60597 => X"89",  -- 137
        60598 => X"80",  -- 128
        60599 => X"6D",  -- 109
        60600 => X"54",  -- 84
        60601 => X"76",  -- 118
        60602 => X"83",  -- 131
        60603 => X"67",  -- 103
        60604 => X"50",  -- 80
        60605 => X"61",  -- 97
        60606 => X"84",  -- 132
        60607 => X"99",  -- 153
        60608 => X"85",  -- 133
        60609 => X"74",  -- 116
        60610 => X"64",  -- 100
        60611 => X"69",  -- 105
        60612 => X"57",  -- 87
        60613 => X"3C",  -- 60
        60614 => X"3C",  -- 60
        60615 => X"7D",  -- 125
        60616 => X"A1",  -- 161
        60617 => X"A9",  -- 169
        60618 => X"85",  -- 133
        60619 => X"2A",  -- 42
        60620 => X"2E",  -- 46
        60621 => X"3C",  -- 60
        60622 => X"90",  -- 144
        60623 => X"7F",  -- 127
        60624 => X"35",  -- 53
        60625 => X"80",  -- 128
        60626 => X"70",  -- 112
        60627 => X"25",  -- 37
        60628 => X"70",  -- 112
        60629 => X"81",  -- 129
        60630 => X"29",  -- 41
        60631 => X"8A",  -- 138
        60632 => X"51",  -- 81
        60633 => X"3B",  -- 59
        60634 => X"31",  -- 49
        60635 => X"3C",  -- 60
        60636 => X"42",  -- 66
        60637 => X"38",  -- 56
        60638 => X"2F",  -- 47
        60639 => X"32",  -- 50
        60640 => X"3C",  -- 60
        60641 => X"37",  -- 55
        60642 => X"3C",  -- 60
        60643 => X"31",  -- 49
        60644 => X"4B",  -- 75
        60645 => X"5C",  -- 92
        60646 => X"2A",  -- 42
        60647 => X"16",  -- 22
        60648 => X"14",  -- 20
        60649 => X"22",  -- 34
        60650 => X"38",  -- 56
        60651 => X"2C",  -- 44
        60652 => X"2F",  -- 47
        60653 => X"27",  -- 39
        60654 => X"27",  -- 39
        60655 => X"32",  -- 50
        60656 => X"2F",  -- 47
        60657 => X"36",  -- 54
        60658 => X"37",  -- 55
        60659 => X"2F",  -- 47
        60660 => X"28",  -- 40
        60661 => X"2B",  -- 43
        60662 => X"33",  -- 51
        60663 => X"3A",  -- 58
        60664 => X"3F",  -- 63
        60665 => X"40",  -- 64
        60666 => X"44",  -- 68
        60667 => X"44",  -- 68
        60668 => X"3E",  -- 62
        60669 => X"39",  -- 57
        60670 => X"3E",  -- 62
        60671 => X"48",  -- 72
        60672 => X"5F",  -- 95
        60673 => X"6D",  -- 109
        60674 => X"75",  -- 117
        60675 => X"6B",  -- 107
        60676 => X"63",  -- 99
        60677 => X"5E",  -- 94
        60678 => X"59",  -- 89
        60679 => X"4F",  -- 79
        60680 => X"4E",  -- 78
        60681 => X"48",  -- 72
        60682 => X"3D",  -- 61
        60683 => X"31",  -- 49
        60684 => X"2A",  -- 42
        60685 => X"28",  -- 40
        60686 => X"29",  -- 41
        60687 => X"29",  -- 41
        60688 => X"2C",  -- 44
        60689 => X"2C",  -- 44
        60690 => X"31",  -- 49
        60691 => X"57",  -- 87
        60692 => X"7A",  -- 122
        60693 => X"8C",  -- 140
        60694 => X"99",  -- 153
        60695 => X"97",  -- 151
        60696 => X"97",  -- 151
        60697 => X"98",  -- 152
        60698 => X"95",  -- 149
        60699 => X"9E",  -- 158
        60700 => X"AD",  -- 173
        60701 => X"9E",  -- 158
        60702 => X"8C",  -- 140
        60703 => X"8F",  -- 143
        60704 => X"87",  -- 135
        60705 => X"8A",  -- 138
        60706 => X"7E",  -- 126
        60707 => X"85",  -- 133
        60708 => X"8D",  -- 141
        60709 => X"84",  -- 132
        60710 => X"8E",  -- 142
        60711 => X"A6",  -- 166
        60712 => X"BB",  -- 187
        60713 => X"BD",  -- 189
        60714 => X"B1",  -- 177
        60715 => X"B5",  -- 181
        60716 => X"B5",  -- 181
        60717 => X"9F",  -- 159
        60718 => X"5A",  -- 90
        60719 => X"32",  -- 50
        60720 => X"96",  -- 150
        60721 => X"9D",  -- 157
        60722 => X"87",  -- 135
        60723 => X"A4",  -- 164
        60724 => X"B4",  -- 180
        60725 => X"9B",  -- 155
        60726 => X"A1",  -- 161
        60727 => X"C0",  -- 192
        60728 => X"C7",  -- 199
        60729 => X"C1",  -- 193
        60730 => X"C6",  -- 198
        60731 => X"D3",  -- 211
        60732 => X"D8",  -- 216
        60733 => X"D1",  -- 209
        60734 => X"CE",  -- 206
        60735 => X"D0",  -- 208
        60736 => X"D4",  -- 212
        60737 => X"DE",  -- 222
        60738 => X"D3",  -- 211
        60739 => X"8C",  -- 140
        60740 => X"80",  -- 128
        60741 => X"B9",  -- 185
        60742 => X"CA",  -- 202
        60743 => X"C5",  -- 197
        60744 => X"D3",  -- 211
        60745 => X"C7",  -- 199
        60746 => X"C4",  -- 196
        60747 => X"C4",  -- 196
        60748 => X"C0",  -- 192
        60749 => X"C3",  -- 195
        60750 => X"CC",  -- 204
        60751 => X"CE",  -- 206
        60752 => X"CE",  -- 206
        60753 => X"D6",  -- 214
        60754 => X"CA",  -- 202
        60755 => X"E4",  -- 228
        60756 => X"97",  -- 151
        60757 => X"2D",  -- 45
        60758 => X"2F",  -- 47
        60759 => X"34",  -- 52
        60760 => X"33",  -- 51
        60761 => X"31",  -- 49
        60762 => X"2C",  -- 44
        60763 => X"2D",  -- 45
        60764 => X"30",  -- 48
        60765 => X"28",  -- 40
        60766 => X"25",  -- 37
        60767 => X"2D",  -- 45
        60768 => X"2A",  -- 42
        60769 => X"25",  -- 37
        60770 => X"25",  -- 37
        60771 => X"28",  -- 40
        60772 => X"25",  -- 37
        60773 => X"1F",  -- 31
        60774 => X"1E",  -- 30
        60775 => X"24",  -- 36
        60776 => X"21",  -- 33
        60777 => X"23",  -- 35
        60778 => X"24",  -- 36
        60779 => X"23",  -- 35
        60780 => X"27",  -- 39
        60781 => X"32",  -- 50
        60782 => X"3E",  -- 62
        60783 => X"44",  -- 68
        60784 => X"45",  -- 69
        60785 => X"54",  -- 84
        60786 => X"60",  -- 96
        60787 => X"63",  -- 99
        60788 => X"69",  -- 105
        60789 => X"74",  -- 116
        60790 => X"7A",  -- 122
        60791 => X"76",  -- 118
        60792 => X"7B",  -- 123
        60793 => X"82",  -- 130
        60794 => X"80",  -- 128
        60795 => X"7E",  -- 126
        60796 => X"83",  -- 131
        60797 => X"82",  -- 130
        60798 => X"82",  -- 130
        60799 => X"8A",  -- 138
        60800 => X"61",  -- 97
        60801 => X"65",  -- 101
        60802 => X"67",  -- 103
        60803 => X"64",  -- 100
        60804 => X"64",  -- 100
        60805 => X"69",  -- 105
        60806 => X"6E",  -- 110
        60807 => X"6E",  -- 110
        60808 => X"6E",  -- 110
        60809 => X"6E",  -- 110
        60810 => X"6F",  -- 111
        60811 => X"70",  -- 112
        60812 => X"72",  -- 114
        60813 => X"73",  -- 115
        60814 => X"71",  -- 113
        60815 => X"6E",  -- 110
        60816 => X"65",  -- 101
        60817 => X"60",  -- 96
        60818 => X"5E",  -- 94
        60819 => X"63",  -- 99
        60820 => X"65",  -- 101
        60821 => X"62",  -- 98
        60822 => X"5D",  -- 93
        60823 => X"5B",  -- 91
        60824 => X"50",  -- 80
        60825 => X"8A",  -- 138
        60826 => X"66",  -- 102
        60827 => X"57",  -- 87
        60828 => X"78",  -- 120
        60829 => X"5F",  -- 95
        60830 => X"56",  -- 86
        60831 => X"83",  -- 131
        60832 => X"7A",  -- 122
        60833 => X"5F",  -- 95
        60834 => X"74",  -- 116
        60835 => X"A0",  -- 160
        60836 => X"72",  -- 114
        60837 => X"58",  -- 88
        60838 => X"9C",  -- 156
        60839 => X"B2",  -- 178
        60840 => X"6B",  -- 107
        60841 => X"53",  -- 83
        60842 => X"44",  -- 68
        60843 => X"4D",  -- 77
        60844 => X"48",  -- 72
        60845 => X"5D",  -- 93
        60846 => X"6D",  -- 109
        60847 => X"3E",  -- 62
        60848 => X"26",  -- 38
        60849 => X"73",  -- 115
        60850 => X"7A",  -- 122
        60851 => X"33",  -- 51
        60852 => X"35",  -- 53
        60853 => X"34",  -- 52
        60854 => X"54",  -- 84
        60855 => X"45",  -- 69
        60856 => X"4E",  -- 78
        60857 => X"93",  -- 147
        60858 => X"64",  -- 100
        60859 => X"25",  -- 37
        60860 => X"26",  -- 38
        60861 => X"74",  -- 116
        60862 => X"88",  -- 136
        60863 => X"3D",  -- 61
        60864 => X"52",  -- 82
        60865 => X"3E",  -- 62
        60866 => X"30",  -- 48
        60867 => X"43",  -- 67
        60868 => X"60",  -- 96
        60869 => X"60",  -- 96
        60870 => X"61",  -- 97
        60871 => X"80",  -- 128
        60872 => X"7A",  -- 122
        60873 => X"64",  -- 100
        60874 => X"63",  -- 99
        60875 => X"72",  -- 114
        60876 => X"84",  -- 132
        60877 => X"61",  -- 97
        60878 => X"59",  -- 89
        60879 => X"6C",  -- 108
        60880 => X"6F",  -- 111
        60881 => X"63",  -- 99
        60882 => X"64",  -- 100
        60883 => X"5E",  -- 94
        60884 => X"6A",  -- 106
        60885 => X"6B",  -- 107
        60886 => X"70",  -- 112
        60887 => X"62",  -- 98
        60888 => X"4D",  -- 77
        60889 => X"33",  -- 51
        60890 => X"13",  -- 19
        60891 => X"02",  -- 2
        60892 => X"03",  -- 3
        60893 => X"07",  -- 7
        60894 => X"07",  -- 7
        60895 => X"08",  -- 8
        60896 => X"0E",  -- 14
        60897 => X"3C",  -- 60
        60898 => X"4A",  -- 74
        60899 => X"71",  -- 113
        60900 => X"6D",  -- 109
        60901 => X"6D",  -- 109
        60902 => X"76",  -- 118
        60903 => X"6F",  -- 111
        60904 => X"7A",  -- 122
        60905 => X"7C",  -- 124
        60906 => X"89",  -- 137
        60907 => X"7A",  -- 122
        60908 => X"6C",  -- 108
        60909 => X"69",  -- 105
        60910 => X"68",  -- 104
        60911 => X"86",  -- 134
        60912 => X"85",  -- 133
        60913 => X"7E",  -- 126
        60914 => X"87",  -- 135
        60915 => X"8F",  -- 143
        60916 => X"A0",  -- 160
        60917 => X"A5",  -- 165
        60918 => X"76",  -- 118
        60919 => X"42",  -- 66
        60920 => X"1E",  -- 30
        60921 => X"1F",  -- 31
        60922 => X"48",  -- 72
        60923 => X"75",  -- 117
        60924 => X"6F",  -- 111
        60925 => X"5A",  -- 90
        60926 => X"5E",  -- 94
        60927 => X"6C",  -- 108
        60928 => X"9F",  -- 159
        60929 => X"A2",  -- 162
        60930 => X"68",  -- 104
        60931 => X"82",  -- 130
        60932 => X"8A",  -- 138
        60933 => X"34",  -- 52
        60934 => X"39",  -- 57
        60935 => X"3E",  -- 62
        60936 => X"53",  -- 83
        60937 => X"91",  -- 145
        60938 => X"DA",  -- 218
        60939 => X"AB",  -- 171
        60940 => X"35",  -- 53
        60941 => X"2A",  -- 42
        60942 => X"3C",  -- 60
        60943 => X"5C",  -- 92
        60944 => X"A4",  -- 164
        60945 => X"67",  -- 103
        60946 => X"64",  -- 100
        60947 => X"74",  -- 116
        60948 => X"39",  -- 57
        60949 => X"50",  -- 80
        60950 => X"87",  -- 135
        60951 => X"4A",  -- 74
        60952 => X"7B",  -- 123
        60953 => X"4C",  -- 76
        60954 => X"36",  -- 54
        60955 => X"35",  -- 53
        60956 => X"2E",  -- 46
        60957 => X"37",  -- 55
        60958 => X"43",  -- 67
        60959 => X"3A",  -- 58
        60960 => X"39",  -- 57
        60961 => X"43",  -- 67
        60962 => X"54",  -- 84
        60963 => X"44",  -- 68
        60964 => X"18",  -- 24
        60965 => X"42",  -- 66
        60966 => X"6E",  -- 110
        60967 => X"29",  -- 41
        60968 => X"16",  -- 22
        60969 => X"16",  -- 22
        60970 => X"37",  -- 55
        60971 => X"2B",  -- 43
        60972 => X"24",  -- 36
        60973 => X"19",  -- 25
        60974 => X"1A",  -- 26
        60975 => X"22",  -- 34
        60976 => X"1B",  -- 27
        60977 => X"24",  -- 36
        60978 => X"26",  -- 38
        60979 => X"20",  -- 32
        60980 => X"19",  -- 25
        60981 => X"1E",  -- 30
        60982 => X"2C",  -- 44
        60983 => X"37",  -- 55
        60984 => X"3F",  -- 63
        60985 => X"42",  -- 66
        60986 => X"46",  -- 70
        60987 => X"47",  -- 71
        60988 => X"43",  -- 67
        60989 => X"3D",  -- 61
        60990 => X"3E",  -- 62
        60991 => X"40",  -- 64
        60992 => X"58",  -- 88
        60993 => X"69",  -- 105
        60994 => X"71",  -- 113
        60995 => X"6B",  -- 107
        60996 => X"63",  -- 99
        60997 => X"5D",  -- 93
        60998 => X"52",  -- 82
        60999 => X"43",  -- 67
        61000 => X"3B",  -- 59
        61001 => X"34",  -- 52
        61002 => X"2C",  -- 44
        61003 => X"24",  -- 36
        61004 => X"21",  -- 33
        61005 => X"21",  -- 33
        61006 => X"24",  -- 36
        61007 => X"26",  -- 38
        61008 => X"2B",  -- 43
        61009 => X"30",  -- 48
        61010 => X"37",  -- 55
        61011 => X"64",  -- 100
        61012 => X"86",  -- 134
        61013 => X"8F",  -- 143
        61014 => X"9C",  -- 156
        61015 => X"96",  -- 150
        61016 => X"90",  -- 144
        61017 => X"96",  -- 150
        61018 => X"98",  -- 152
        61019 => X"9C",  -- 156
        61020 => X"A3",  -- 163
        61021 => X"9C",  -- 156
        61022 => X"94",  -- 148
        61023 => X"95",  -- 149
        61024 => X"91",  -- 145
        61025 => X"79",  -- 121
        61026 => X"72",  -- 114
        61027 => X"72",  -- 114
        61028 => X"78",  -- 120
        61029 => X"84",  -- 132
        61030 => X"8B",  -- 139
        61031 => X"96",  -- 150
        61032 => X"B4",  -- 180
        61033 => X"B9",  -- 185
        61034 => X"B6",  -- 182
        61035 => X"B3",  -- 179
        61036 => X"B1",  -- 177
        61037 => X"8C",  -- 140
        61038 => X"2D",  -- 45
        61039 => X"24",  -- 36
        61040 => X"81",  -- 129
        61041 => X"A3",  -- 163
        61042 => X"8A",  -- 138
        61043 => X"A9",  -- 169
        61044 => X"B0",  -- 176
        61045 => X"A5",  -- 165
        61046 => X"A7",  -- 167
        61047 => X"C0",  -- 192
        61048 => X"CA",  -- 202
        61049 => X"C7",  -- 199
        61050 => X"C8",  -- 200
        61051 => X"CA",  -- 202
        61052 => X"CD",  -- 205
        61053 => X"CF",  -- 207
        61054 => X"CE",  -- 206
        61055 => X"CE",  -- 206
        61056 => X"D6",  -- 214
        61057 => X"DB",  -- 219
        61058 => X"DF",  -- 223
        61059 => X"A3",  -- 163
        61060 => X"84",  -- 132
        61061 => X"AF",  -- 175
        61062 => X"C9",  -- 201
        61063 => X"CF",  -- 207
        61064 => X"D5",  -- 213
        61065 => X"CC",  -- 204
        61066 => X"CD",  -- 205
        61067 => X"CD",  -- 205
        61068 => X"C8",  -- 200
        61069 => X"CA",  -- 202
        61070 => X"D1",  -- 209
        61071 => X"D1",  -- 209
        61072 => X"CE",  -- 206
        61073 => X"DB",  -- 219
        61074 => X"D2",  -- 210
        61075 => X"E1",  -- 225
        61076 => X"BB",  -- 187
        61077 => X"4B",  -- 75
        61078 => X"2E",  -- 46
        61079 => X"36",  -- 54
        61080 => X"37",  -- 55
        61081 => X"32",  -- 50
        61082 => X"2A",  -- 42
        61083 => X"2A",  -- 42
        61084 => X"2F",  -- 47
        61085 => X"29",  -- 41
        61086 => X"24",  -- 36
        61087 => X"2D",  -- 45
        61088 => X"2B",  -- 43
        61089 => X"27",  -- 39
        61090 => X"28",  -- 40
        61091 => X"2C",  -- 44
        61092 => X"29",  -- 41
        61093 => X"20",  -- 32
        61094 => X"1F",  -- 31
        61095 => X"24",  -- 36
        61096 => X"23",  -- 35
        61097 => X"28",  -- 40
        61098 => X"2B",  -- 43
        61099 => X"2A",  -- 42
        61100 => X"2D",  -- 45
        61101 => X"38",  -- 56
        61102 => X"42",  -- 66
        61103 => X"48",  -- 72
        61104 => X"4E",  -- 78
        61105 => X"5F",  -- 95
        61106 => X"68",  -- 104
        61107 => X"65",  -- 101
        61108 => X"66",  -- 102
        61109 => X"72",  -- 114
        61110 => X"79",  -- 121
        61111 => X"78",  -- 120
        61112 => X"81",  -- 129
        61113 => X"85",  -- 133
        61114 => X"7F",  -- 127
        61115 => X"7B",  -- 123
        61116 => X"7F",  -- 127
        61117 => X"7E",  -- 126
        61118 => X"80",  -- 128
        61119 => X"88",  -- 136
        61120 => X"61",  -- 97
        61121 => X"63",  -- 99
        61122 => X"61",  -- 97
        61123 => X"5D",  -- 93
        61124 => X"5D",  -- 93
        61125 => X"5F",  -- 95
        61126 => X"60",  -- 96
        61127 => X"5C",  -- 92
        61128 => X"6E",  -- 110
        61129 => X"6E",  -- 110
        61130 => X"71",  -- 113
        61131 => X"6E",  -- 110
        61132 => X"6C",  -- 108
        61133 => X"69",  -- 105
        61134 => X"68",  -- 104
        61135 => X"68",  -- 104
        61136 => X"63",  -- 99
        61137 => X"61",  -- 97
        61138 => X"64",  -- 100
        61139 => X"6C",  -- 108
        61140 => X"6D",  -- 109
        61141 => X"67",  -- 103
        61142 => X"69",  -- 105
        61143 => X"71",  -- 113
        61144 => X"89",  -- 137
        61145 => X"5A",  -- 90
        61146 => X"5C",  -- 92
        61147 => X"5F",  -- 95
        61148 => X"49",  -- 73
        61149 => X"5C",  -- 92
        61150 => X"7F",  -- 127
        61151 => X"81",  -- 129
        61152 => X"5D",  -- 93
        61153 => X"8A",  -- 138
        61154 => X"94",  -- 148
        61155 => X"64",  -- 100
        61156 => X"4A",  -- 74
        61157 => X"81",  -- 129
        61158 => X"A7",  -- 167
        61159 => X"64",  -- 100
        61160 => X"66",  -- 102
        61161 => X"6C",  -- 108
        61162 => X"72",  -- 114
        61163 => X"60",  -- 96
        61164 => X"68",  -- 104
        61165 => X"7F",  -- 127
        61166 => X"70",  -- 112
        61167 => X"5A",  -- 90
        61168 => X"75",  -- 117
        61169 => X"7C",  -- 124
        61170 => X"4A",  -- 74
        61171 => X"22",  -- 34
        61172 => X"37",  -- 55
        61173 => X"63",  -- 99
        61174 => X"58",  -- 88
        61175 => X"57",  -- 87
        61176 => X"9A",  -- 154
        61177 => X"7E",  -- 126
        61178 => X"34",  -- 52
        61179 => X"25",  -- 37
        61180 => X"7F",  -- 127
        61181 => X"81",  -- 129
        61182 => X"37",  -- 55
        61183 => X"69",  -- 105
        61184 => X"67",  -- 103
        61185 => X"48",  -- 72
        61186 => X"3C",  -- 60
        61187 => X"4A",  -- 74
        61188 => X"2E",  -- 46
        61189 => X"1F",  -- 31
        61190 => X"4A",  -- 74
        61191 => X"55",  -- 85
        61192 => X"39",  -- 57
        61193 => X"4B",  -- 75
        61194 => X"63",  -- 99
        61195 => X"6B",  -- 107
        61196 => X"77",  -- 119
        61197 => X"58",  -- 88
        61198 => X"51",  -- 81
        61199 => X"5F",  -- 95
        61200 => X"5F",  -- 95
        61201 => X"6F",  -- 111
        61202 => X"67",  -- 103
        61203 => X"51",  -- 81
        61204 => X"65",  -- 101
        61205 => X"56",  -- 86
        61206 => X"48",  -- 72
        61207 => X"49",  -- 73
        61208 => X"24",  -- 36
        61209 => X"15",  -- 21
        61210 => X"10",  -- 16
        61211 => X"14",  -- 20
        61212 => X"12",  -- 18
        61213 => X"12",  -- 18
        61214 => X"12",  -- 18
        61215 => X"0C",  -- 12
        61216 => X"09",  -- 9
        61217 => X"2B",  -- 43
        61218 => X"39",  -- 57
        61219 => X"48",  -- 72
        61220 => X"63",  -- 99
        61221 => X"5F",  -- 95
        61222 => X"80",  -- 128
        61223 => X"68",  -- 104
        61224 => X"5F",  -- 95
        61225 => X"64",  -- 100
        61226 => X"7E",  -- 126
        61227 => X"6C",  -- 108
        61228 => X"63",  -- 99
        61229 => X"6C",  -- 108
        61230 => X"68",  -- 104
        61231 => X"91",  -- 145
        61232 => X"7E",  -- 126
        61233 => X"77",  -- 119
        61234 => X"76",  -- 118
        61235 => X"57",  -- 87
        61236 => X"59",  -- 89
        61237 => X"73",  -- 115
        61238 => X"4F",  -- 79
        61239 => X"21",  -- 33
        61240 => X"25",  -- 37
        61241 => X"25",  -- 37
        61242 => X"50",  -- 80
        61243 => X"7E",  -- 126
        61244 => X"7E",  -- 126
        61245 => X"71",  -- 113
        61246 => X"67",  -- 103
        61247 => X"55",  -- 85
        61248 => X"73",  -- 115
        61249 => X"78",  -- 120
        61250 => X"8F",  -- 143
        61251 => X"80",  -- 128
        61252 => X"8A",  -- 138
        61253 => X"4B",  -- 75
        61254 => X"3B",  -- 59
        61255 => X"43",  -- 67
        61256 => X"3F",  -- 63
        61257 => X"38",  -- 56
        61258 => X"6B",  -- 107
        61259 => X"D5",  -- 213
        61260 => X"A1",  -- 161
        61261 => X"3E",  -- 62
        61262 => X"39",  -- 57
        61263 => X"3A",  -- 58
        61264 => X"43",  -- 67
        61265 => X"70",  -- 112
        61266 => X"8A",  -- 138
        61267 => X"79",  -- 121
        61268 => X"73",  -- 115
        61269 => X"3F",  -- 63
        61270 => X"67",  -- 103
        61271 => X"88",  -- 136
        61272 => X"56",  -- 86
        61273 => X"6B",  -- 107
        61274 => X"52",  -- 82
        61275 => X"32",  -- 50
        61276 => X"3A",  -- 58
        61277 => X"39",  -- 57
        61278 => X"2F",  -- 47
        61279 => X"3D",  -- 61
        61280 => X"3D",  -- 61
        61281 => X"49",  -- 73
        61282 => X"3F",  -- 63
        61283 => X"38",  -- 56
        61284 => X"34",  -- 52
        61285 => X"0A",  -- 10
        61286 => X"18",  -- 24
        61287 => X"7E",  -- 126
        61288 => X"3C",  -- 60
        61289 => X"17",  -- 23
        61290 => X"21",  -- 33
        61291 => X"14",  -- 20
        61292 => X"17",  -- 23
        61293 => X"16",  -- 22
        61294 => X"15",  -- 21
        61295 => X"12",  -- 18
        61296 => X"10",  -- 16
        61297 => X"14",  -- 20
        61298 => X"14",  -- 20
        61299 => X"13",  -- 19
        61300 => X"18",  -- 24
        61301 => X"24",  -- 36
        61302 => X"32",  -- 50
        61303 => X"39",  -- 57
        61304 => X"36",  -- 54
        61305 => X"38",  -- 56
        61306 => X"3E",  -- 62
        61307 => X"45",  -- 69
        61308 => X"48",  -- 72
        61309 => X"46",  -- 70
        61310 => X"43",  -- 67
        61311 => X"43",  -- 67
        61312 => X"50",  -- 80
        61313 => X"61",  -- 97
        61314 => X"69",  -- 105
        61315 => X"65",  -- 101
        61316 => X"5F",  -- 95
        61317 => X"58",  -- 88
        61318 => X"49",  -- 73
        61319 => X"36",  -- 54
        61320 => X"30",  -- 48
        61321 => X"2A",  -- 42
        61322 => X"25",  -- 37
        61323 => X"22",  -- 34
        61324 => X"23",  -- 35
        61325 => X"25",  -- 37
        61326 => X"28",  -- 40
        61327 => X"2A",  -- 42
        61328 => X"2F",  -- 47
        61329 => X"39",  -- 57
        61330 => X"42",  -- 66
        61331 => X"70",  -- 112
        61332 => X"91",  -- 145
        61333 => X"97",  -- 151
        61334 => X"A3",  -- 163
        61335 => X"9C",  -- 156
        61336 => X"8F",  -- 143
        61337 => X"95",  -- 149
        61338 => X"96",  -- 150
        61339 => X"91",  -- 145
        61340 => X"91",  -- 145
        61341 => X"95",  -- 149
        61342 => X"94",  -- 148
        61343 => X"8F",  -- 143
        61344 => X"75",  -- 117
        61345 => X"4E",  -- 78
        61346 => X"5F",  -- 95
        61347 => X"6D",  -- 109
        61348 => X"78",  -- 120
        61349 => X"99",  -- 153
        61350 => X"A0",  -- 160
        61351 => X"97",  -- 151
        61352 => X"A8",  -- 168
        61353 => X"A6",  -- 166
        61354 => X"AB",  -- 171
        61355 => X"B2",  -- 178
        61356 => X"AA",  -- 170
        61357 => X"70",  -- 112
        61358 => X"05",  -- 5
        61359 => X"24",  -- 36
        61360 => X"61",  -- 97
        61361 => X"9F",  -- 159
        61362 => X"81",  -- 129
        61363 => X"96",  -- 150
        61364 => X"A1",  -- 161
        61365 => X"B6",  -- 182
        61366 => X"B1",  -- 177
        61367 => X"AE",  -- 174
        61368 => X"C6",  -- 198
        61369 => X"CC",  -- 204
        61370 => X"CC",  -- 204
        61371 => X"C9",  -- 201
        61372 => X"CB",  -- 203
        61373 => X"D3",  -- 211
        61374 => X"D6",  -- 214
        61375 => X"D2",  -- 210
        61376 => X"D4",  -- 212
        61377 => X"D4",  -- 212
        61378 => X"E9",  -- 233
        61379 => X"BF",  -- 191
        61380 => X"90",  -- 144
        61381 => X"A6",  -- 166
        61382 => X"C0",  -- 192
        61383 => X"D3",  -- 211
        61384 => X"D4",  -- 212
        61385 => X"CE",  -- 206
        61386 => X"D5",  -- 213
        61387 => X"DB",  -- 219
        61388 => X"D8",  -- 216
        61389 => X"D6",  -- 214
        61390 => X"D8",  -- 216
        61391 => X"D4",  -- 212
        61392 => X"D6",  -- 214
        61393 => X"DA",  -- 218
        61394 => X"D3",  -- 211
        61395 => X"D3",  -- 211
        61396 => X"CF",  -- 207
        61397 => X"6A",  -- 106
        61398 => X"32",  -- 50
        61399 => X"39",  -- 57
        61400 => X"39",  -- 57
        61401 => X"31",  -- 49
        61402 => X"28",  -- 40
        61403 => X"28",  -- 40
        61404 => X"2F",  -- 47
        61405 => X"29",  -- 41
        61406 => X"25",  -- 37
        61407 => X"2C",  -- 44
        61408 => X"2C",  -- 44
        61409 => X"28",  -- 40
        61410 => X"2A",  -- 42
        61411 => X"2E",  -- 46
        61412 => X"2D",  -- 45
        61413 => X"23",  -- 35
        61414 => X"20",  -- 32
        61415 => X"22",  -- 34
        61416 => X"27",  -- 39
        61417 => X"2D",  -- 45
        61418 => X"32",  -- 50
        61419 => X"31",  -- 49
        61420 => X"35",  -- 53
        61421 => X"3D",  -- 61
        61422 => X"48",  -- 72
        61423 => X"4A",  -- 74
        61424 => X"56",  -- 86
        61425 => X"66",  -- 102
        61426 => X"6D",  -- 109
        61427 => X"66",  -- 102
        61428 => X"63",  -- 99
        61429 => X"6F",  -- 111
        61430 => X"7B",  -- 123
        61431 => X"7D",  -- 125
        61432 => X"87",  -- 135
        61433 => X"88",  -- 136
        61434 => X"7F",  -- 127
        61435 => X"79",  -- 121
        61436 => X"7B",  -- 123
        61437 => X"7B",  -- 123
        61438 => X"7E",  -- 126
        61439 => X"87",  -- 135
        61440 => X"4D",  -- 77
        61441 => X"50",  -- 80
        61442 => X"55",  -- 85
        61443 => X"58",  -- 88
        61444 => X"5A",  -- 90
        61445 => X"5C",  -- 92
        61446 => X"5D",  -- 93
        61447 => X"5F",  -- 95
        61448 => X"65",  -- 101
        61449 => X"67",  -- 103
        61450 => X"69",  -- 105
        61451 => X"6A",  -- 106
        61452 => X"6F",  -- 111
        61453 => X"6F",  -- 111
        61454 => X"65",  -- 101
        61455 => X"58",  -- 88
        61456 => X"4E",  -- 78
        61457 => X"61",  -- 97
        61458 => X"69",  -- 105
        61459 => X"5E",  -- 94
        61460 => X"5F",  -- 95
        61461 => X"79",  -- 121
        61462 => X"86",  -- 134
        61463 => X"78",  -- 120
        61464 => X"61",  -- 97
        61465 => X"52",  -- 82
        61466 => X"51",  -- 81
        61467 => X"54",  -- 84
        61468 => X"5B",  -- 91
        61469 => X"71",  -- 113
        61470 => X"7A",  -- 122
        61471 => X"6D",  -- 109
        61472 => X"94",  -- 148
        61473 => X"79",  -- 121
        61474 => X"6B",  -- 107
        61475 => X"5C",  -- 92
        61476 => X"9F",  -- 159
        61477 => X"B0",  -- 176
        61478 => X"56",  -- 86
        61479 => X"5C",  -- 92
        61480 => X"69",  -- 105
        61481 => X"69",  -- 105
        61482 => X"66",  -- 102
        61483 => X"5D",  -- 93
        61484 => X"76",  -- 118
        61485 => X"79",  -- 121
        61486 => X"61",  -- 97
        61487 => X"87",  -- 135
        61488 => X"81",  -- 129
        61489 => X"5E",  -- 94
        61490 => X"44",  -- 68
        61491 => X"45",  -- 69
        61492 => X"75",  -- 117
        61493 => X"5E",  -- 94
        61494 => X"62",  -- 98
        61495 => X"A6",  -- 166
        61496 => X"85",  -- 133
        61497 => X"5E",  -- 94
        61498 => X"3D",  -- 61
        61499 => X"72",  -- 114
        61500 => X"82",  -- 130
        61501 => X"3D",  -- 61
        61502 => X"60",  -- 96
        61503 => X"83",  -- 131
        61504 => X"63",  -- 99
        61505 => X"5E",  -- 94
        61506 => X"75",  -- 117
        61507 => X"42",  -- 66
        61508 => X"35",  -- 53
        61509 => X"1D",  -- 29
        61510 => X"39",  -- 57
        61511 => X"23",  -- 35
        61512 => X"29",  -- 41
        61513 => X"0C",  -- 12
        61514 => X"33",  -- 51
        61515 => X"44",  -- 68
        61516 => X"36",  -- 54
        61517 => X"3C",  -- 60
        61518 => X"41",  -- 65
        61519 => X"62",  -- 98
        61520 => X"6F",  -- 111
        61521 => X"60",  -- 96
        61522 => X"64",  -- 100
        61523 => X"63",  -- 99
        61524 => X"54",  -- 84
        61525 => X"3B",  -- 59
        61526 => X"1F",  -- 31
        61527 => X"20",  -- 32
        61528 => X"1C",  -- 28
        61529 => X"11",  -- 17
        61530 => X"11",  -- 17
        61531 => X"21",  -- 33
        61532 => X"32",  -- 50
        61533 => X"3F",  -- 63
        61534 => X"3A",  -- 58
        61535 => X"29",  -- 41
        61536 => X"43",  -- 67
        61537 => X"39",  -- 57
        61538 => X"29",  -- 41
        61539 => X"32",  -- 50
        61540 => X"3A",  -- 58
        61541 => X"49",  -- 73
        61542 => X"72",  -- 114
        61543 => X"65",  -- 101
        61544 => X"61",  -- 97
        61545 => X"75",  -- 117
        61546 => X"66",  -- 102
        61547 => X"6F",  -- 111
        61548 => X"60",  -- 96
        61549 => X"5E",  -- 94
        61550 => X"5B",  -- 91
        61551 => X"4D",  -- 77
        61552 => X"63",  -- 99
        61553 => X"6C",  -- 108
        61554 => X"27",  -- 39
        61555 => X"13",  -- 19
        61556 => X"1D",  -- 29
        61557 => X"5B",  -- 91
        61558 => X"2A",  -- 42
        61559 => X"3E",  -- 62
        61560 => X"39",  -- 57
        61561 => X"45",  -- 69
        61562 => X"53",  -- 83
        61563 => X"44",  -- 68
        61564 => X"7A",  -- 122
        61565 => X"80",  -- 128
        61566 => X"67",  -- 103
        61567 => X"75",  -- 117
        61568 => X"76",  -- 118
        61569 => X"78",  -- 120
        61570 => X"66",  -- 102
        61571 => X"9B",  -- 155
        61572 => X"8D",  -- 141
        61573 => X"7F",  -- 127
        61574 => X"4B",  -- 75
        61575 => X"39",  -- 57
        61576 => X"43",  -- 67
        61577 => X"41",  -- 65
        61578 => X"32",  -- 50
        61579 => X"49",  -- 73
        61580 => X"C1",  -- 193
        61581 => X"88",  -- 136
        61582 => X"31",  -- 49
        61583 => X"43",  -- 67
        61584 => X"44",  -- 68
        61585 => X"41",  -- 65
        61586 => X"4F",  -- 79
        61587 => X"8F",  -- 143
        61588 => X"79",  -- 121
        61589 => X"83",  -- 131
        61590 => X"4A",  -- 74
        61591 => X"5D",  -- 93
        61592 => X"8E",  -- 142
        61593 => X"4E",  -- 78
        61594 => X"7F",  -- 127
        61595 => X"44",  -- 68
        61596 => X"39",  -- 57
        61597 => X"2E",  -- 46
        61598 => X"3E",  -- 62
        61599 => X"39",  -- 57
        61600 => X"3E",  -- 62
        61601 => X"47",  -- 71
        61602 => X"45",  -- 69
        61603 => X"2F",  -- 47
        61604 => X"19",  -- 25
        61605 => X"11",  -- 17
        61606 => X"0F",  -- 15
        61607 => X"0E",  -- 14
        61608 => X"6D",  -- 109
        61609 => X"5D",  -- 93
        61610 => X"1C",  -- 28
        61611 => X"0C",  -- 12
        61612 => X"15",  -- 21
        61613 => X"13",  -- 19
        61614 => X"0F",  -- 15
        61615 => X"14",  -- 20
        61616 => X"0F",  -- 15
        61617 => X"11",  -- 17
        61618 => X"0F",  -- 15
        61619 => X"0E",  -- 14
        61620 => X"1B",  -- 27
        61621 => X"2D",  -- 45
        61622 => X"38",  -- 56
        61623 => X"37",  -- 55
        61624 => X"3A",  -- 58
        61625 => X"2F",  -- 47
        61626 => X"2B",  -- 43
        61627 => X"35",  -- 53
        61628 => X"3E",  -- 62
        61629 => X"44",  -- 68
        61630 => X"43",  -- 67
        61631 => X"45",  -- 69
        61632 => X"46",  -- 70
        61633 => X"54",  -- 84
        61634 => X"64",  -- 100
        61635 => X"6A",  -- 106
        61636 => X"62",  -- 98
        61637 => X"51",  -- 81
        61638 => X"3C",  -- 60
        61639 => X"2E",  -- 46
        61640 => X"2D",  -- 45
        61641 => X"2F",  -- 47
        61642 => X"2C",  -- 44
        61643 => X"25",  -- 37
        61644 => X"20",  -- 32
        61645 => X"23",  -- 35
        61646 => X"2C",  -- 44
        61647 => X"30",  -- 48
        61648 => X"2D",  -- 45
        61649 => X"42",  -- 66
        61650 => X"47",  -- 71
        61651 => X"81",  -- 129
        61652 => X"87",  -- 135
        61653 => X"98",  -- 152
        61654 => X"B3",  -- 179
        61655 => X"A3",  -- 163
        61656 => X"91",  -- 145
        61657 => X"93",  -- 147
        61658 => X"94",  -- 148
        61659 => X"8D",  -- 141
        61660 => X"94",  -- 148
        61661 => X"94",  -- 148
        61662 => X"85",  -- 133
        61663 => X"8C",  -- 140
        61664 => X"5B",  -- 91
        61665 => X"20",  -- 32
        61666 => X"42",  -- 66
        61667 => X"6C",  -- 108
        61668 => X"8D",  -- 141
        61669 => X"9C",  -- 156
        61670 => X"A5",  -- 165
        61671 => X"A2",  -- 162
        61672 => X"AE",  -- 174
        61673 => X"B2",  -- 178
        61674 => X"9D",  -- 157
        61675 => X"AD",  -- 173
        61676 => X"95",  -- 149
        61677 => X"5D",  -- 93
        61678 => X"05",  -- 5
        61679 => X"1C",  -- 28
        61680 => X"6F",  -- 111
        61681 => X"98",  -- 152
        61682 => X"A1",  -- 161
        61683 => X"79",  -- 121
        61684 => X"7F",  -- 127
        61685 => X"A6",  -- 166
        61686 => X"B4",  -- 180
        61687 => X"B1",  -- 177
        61688 => X"BA",  -- 186
        61689 => X"C5",  -- 197
        61690 => X"C9",  -- 201
        61691 => X"CC",  -- 204
        61692 => X"D6",  -- 214
        61693 => X"DA",  -- 218
        61694 => X"D6",  -- 214
        61695 => X"D8",  -- 216
        61696 => X"DB",  -- 219
        61697 => X"C5",  -- 197
        61698 => X"E6",  -- 230
        61699 => X"D1",  -- 209
        61700 => X"9A",  -- 154
        61701 => X"A7",  -- 167
        61702 => X"C5",  -- 197
        61703 => X"CC",  -- 204
        61704 => X"D5",  -- 213
        61705 => X"D3",  -- 211
        61706 => X"D8",  -- 216
        61707 => X"DD",  -- 221
        61708 => X"DD",  -- 221
        61709 => X"D8",  -- 216
        61710 => X"DA",  -- 218
        61711 => X"E1",  -- 225
        61712 => X"D7",  -- 215
        61713 => X"CF",  -- 207
        61714 => X"D0",  -- 208
        61715 => X"D2",  -- 210
        61716 => X"D0",  -- 208
        61717 => X"92",  -- 146
        61718 => X"3D",  -- 61
        61719 => X"3C",  -- 60
        61720 => X"34",  -- 52
        61721 => X"2D",  -- 45
        61722 => X"2B",  -- 43
        61723 => X"2B",  -- 43
        61724 => X"2A",  -- 42
        61725 => X"27",  -- 39
        61726 => X"26",  -- 38
        61727 => X"28",  -- 40
        61728 => X"27",  -- 39
        61729 => X"29",  -- 41
        61730 => X"2C",  -- 44
        61731 => X"2D",  -- 45
        61732 => X"2C",  -- 44
        61733 => X"29",  -- 41
        61734 => X"25",  -- 37
        61735 => X"22",  -- 34
        61736 => X"2C",  -- 44
        61737 => X"2E",  -- 46
        61738 => X"33",  -- 51
        61739 => X"36",  -- 54
        61740 => X"3C",  -- 60
        61741 => X"44",  -- 68
        61742 => X"50",  -- 80
        61743 => X"57",  -- 87
        61744 => X"59",  -- 89
        61745 => X"66",  -- 102
        61746 => X"6E",  -- 110
        61747 => X"63",  -- 99
        61748 => X"5D",  -- 93
        61749 => X"70",  -- 112
        61750 => X"83",  -- 131
        61751 => X"7F",  -- 127
        61752 => X"82",  -- 130
        61753 => X"8D",  -- 141
        61754 => X"7B",  -- 123
        61755 => X"6A",  -- 106
        61756 => X"75",  -- 117
        61757 => X"76",  -- 118
        61758 => X"72",  -- 114
        61759 => X"82",  -- 130
        61760 => X"4F",  -- 79
        61761 => X"51",  -- 81
        61762 => X"53",  -- 83
        61763 => X"55",  -- 85
        61764 => X"56",  -- 86
        61765 => X"58",  -- 88
        61766 => X"5B",  -- 91
        61767 => X"5E",  -- 94
        61768 => X"51",  -- 81
        61769 => X"53",  -- 83
        61770 => X"55",  -- 85
        61771 => X"5C",  -- 92
        61772 => X"65",  -- 101
        61773 => X"67",  -- 103
        61774 => X"5B",  -- 91
        61775 => X"4D",  -- 77
        61776 => X"56",  -- 86
        61777 => X"5D",  -- 93
        61778 => X"5D",  -- 93
        61779 => X"6D",  -- 109
        61780 => X"88",  -- 136
        61781 => X"7F",  -- 127
        61782 => X"5D",  -- 93
        61783 => X"4C",  -- 76
        61784 => X"5E",  -- 94
        61785 => X"59",  -- 89
        61786 => X"54",  -- 84
        61787 => X"44",  -- 68
        61788 => X"66",  -- 102
        61789 => X"82",  -- 130
        61790 => X"77",  -- 119
        61791 => X"9D",  -- 157
        61792 => X"6D",  -- 109
        61793 => X"5D",  -- 93
        61794 => X"5E",  -- 94
        61795 => X"8A",  -- 138
        61796 => X"91",  -- 145
        61797 => X"6F",  -- 111
        61798 => X"64",  -- 100
        61799 => X"61",  -- 97
        61800 => X"66",  -- 102
        61801 => X"55",  -- 85
        61802 => X"63",  -- 99
        61803 => X"5F",  -- 95
        61804 => X"75",  -- 117
        61805 => X"5D",  -- 93
        61806 => X"6D",  -- 109
        61807 => X"A0",  -- 160
        61808 => X"7A",  -- 122
        61809 => X"51",  -- 81
        61810 => X"54",  -- 84
        61811 => X"76",  -- 118
        61812 => X"6E",  -- 110
        61813 => X"60",  -- 96
        61814 => X"97",  -- 151
        61815 => X"8C",  -- 140
        61816 => X"6D",  -- 109
        61817 => X"45",  -- 69
        61818 => X"7C",  -- 124
        61819 => X"89",  -- 137
        61820 => X"45",  -- 69
        61821 => X"5E",  -- 94
        61822 => X"7B",  -- 123
        61823 => X"7D",  -- 125
        61824 => X"70",  -- 112
        61825 => X"5E",  -- 94
        61826 => X"5A",  -- 90
        61827 => X"47",  -- 71
        61828 => X"43",  -- 67
        61829 => X"57",  -- 87
        61830 => X"37",  -- 55
        61831 => X"3A",  -- 58
        61832 => X"0F",  -- 15
        61833 => X"02",  -- 2
        61834 => X"2C",  -- 44
        61835 => X"2F",  -- 47
        61836 => X"2C",  -- 44
        61837 => X"37",  -- 55
        61838 => X"3F",  -- 63
        61839 => X"55",  -- 85
        61840 => X"53",  -- 83
        61841 => X"4A",  -- 74
        61842 => X"47",  -- 71
        61843 => X"3A",  -- 58
        61844 => X"33",  -- 51
        61845 => X"2F",  -- 47
        61846 => X"19",  -- 25
        61847 => X"10",  -- 16
        61848 => X"26",  -- 38
        61849 => X"22",  -- 34
        61850 => X"23",  -- 35
        61851 => X"38",  -- 56
        61852 => X"54",  -- 84
        61853 => X"59",  -- 89
        61854 => X"3C",  -- 60
        61855 => X"1B",  -- 27
        61856 => X"29",  -- 41
        61857 => X"2E",  -- 46
        61858 => X"27",  -- 39
        61859 => X"26",  -- 38
        61860 => X"15",  -- 21
        61861 => X"20",  -- 32
        61862 => X"4C",  -- 76
        61863 => X"45",  -- 69
        61864 => X"47",  -- 71
        61865 => X"5F",  -- 95
        61866 => X"5D",  -- 93
        61867 => X"54",  -- 84
        61868 => X"5E",  -- 94
        61869 => X"54",  -- 84
        61870 => X"4F",  -- 79
        61871 => X"2F",  -- 47
        61872 => X"27",  -- 39
        61873 => X"52",  -- 82
        61874 => X"55",  -- 85
        61875 => X"14",  -- 20
        61876 => X"1B",  -- 27
        61877 => X"41",  -- 65
        61878 => X"48",  -- 72
        61879 => X"2B",  -- 43
        61880 => X"54",  -- 84
        61881 => X"52",  -- 82
        61882 => X"47",  -- 71
        61883 => X"66",  -- 102
        61884 => X"48",  -- 72
        61885 => X"65",  -- 101
        61886 => X"8E",  -- 142
        61887 => X"60",  -- 96
        61888 => X"74",  -- 116
        61889 => X"6E",  -- 110
        61890 => X"8E",  -- 142
        61891 => X"74",  -- 116
        61892 => X"6F",  -- 111
        61893 => X"94",  -- 148
        61894 => X"A0",  -- 160
        61895 => X"4C",  -- 76
        61896 => X"3C",  -- 60
        61897 => X"46",  -- 70
        61898 => X"47",  -- 71
        61899 => X"3F",  -- 63
        61900 => X"52",  -- 82
        61901 => X"D3",  -- 211
        61902 => X"8B",  -- 139
        61903 => X"3A",  -- 58
        61904 => X"3A",  -- 58
        61905 => X"52",  -- 82
        61906 => X"4C",  -- 76
        61907 => X"48",  -- 72
        61908 => X"85",  -- 133
        61909 => X"79",  -- 121
        61910 => X"84",  -- 132
        61911 => X"52",  -- 82
        61912 => X"58",  -- 88
        61913 => X"81",  -- 129
        61914 => X"58",  -- 88
        61915 => X"6F",  -- 111
        61916 => X"37",  -- 55
        61917 => X"44",  -- 68
        61918 => X"45",  -- 69
        61919 => X"37",  -- 55
        61920 => X"42",  -- 66
        61921 => X"43",  -- 67
        61922 => X"3A",  -- 58
        61923 => X"27",  -- 39
        61924 => X"17",  -- 23
        61925 => X"10",  -- 16
        61926 => X"12",  -- 18
        61927 => X"13",  -- 19
        61928 => X"20",  -- 32
        61929 => X"5B",  -- 91
        61930 => X"59",  -- 89
        61931 => X"1A",  -- 26
        61932 => X"0C",  -- 12
        61933 => X"0C",  -- 12
        61934 => X"1E",  -- 30
        61935 => X"0A",  -- 10
        61936 => X"10",  -- 16
        61937 => X"14",  -- 20
        61938 => X"17",  -- 23
        61939 => X"19",  -- 25
        61940 => X"26",  -- 38
        61941 => X"3A",  -- 58
        61942 => X"44",  -- 68
        61943 => X"45",  -- 69
        61944 => X"34",  -- 52
        61945 => X"2E",  -- 46
        61946 => X"2B",  -- 43
        61947 => X"2F",  -- 47
        61948 => X"32",  -- 50
        61949 => X"33",  -- 51
        61950 => X"34",  -- 52
        61951 => X"39",  -- 57
        61952 => X"46",  -- 70
        61953 => X"52",  -- 82
        61954 => X"62",  -- 98
        61955 => X"6A",  -- 106
        61956 => X"62",  -- 98
        61957 => X"51",  -- 81
        61958 => X"3F",  -- 63
        61959 => X"31",  -- 49
        61960 => X"39",  -- 57
        61961 => X"3A",  -- 58
        61962 => X"39",  -- 57
        61963 => X"2E",  -- 46
        61964 => X"27",  -- 39
        61965 => X"27",  -- 39
        61966 => X"2E",  -- 46
        61967 => X"33",  -- 51
        61968 => X"40",  -- 64
        61969 => X"37",  -- 55
        61970 => X"5D",  -- 93
        61971 => X"92",  -- 146
        61972 => X"92",  -- 146
        61973 => X"98",  -- 152
        61974 => X"9E",  -- 158
        61975 => X"99",  -- 153
        61976 => X"92",  -- 146
        61977 => X"84",  -- 132
        61978 => X"8A",  -- 138
        61979 => X"7D",  -- 125
        61980 => X"75",  -- 117
        61981 => X"8A",  -- 138
        61982 => X"8B",  -- 139
        61983 => X"79",  -- 121
        61984 => X"36",  -- 54
        61985 => X"11",  -- 17
        61986 => X"3A",  -- 58
        61987 => X"90",  -- 144
        61988 => X"9A",  -- 154
        61989 => X"A6",  -- 166
        61990 => X"A0",  -- 160
        61991 => X"BB",  -- 187
        61992 => X"9C",  -- 156
        61993 => X"A1",  -- 161
        61994 => X"A0",  -- 160
        61995 => X"AB",  -- 171
        61996 => X"8E",  -- 142
        61997 => X"2F",  -- 47
        61998 => X"01",  -- 1
        61999 => X"12",  -- 18
        62000 => X"5A",  -- 90
        62001 => X"98",  -- 152
        62002 => X"A5",  -- 165
        62003 => X"78",  -- 120
        62004 => X"81",  -- 129
        62005 => X"B7",  -- 183
        62006 => X"AF",  -- 175
        62007 => X"AC",  -- 172
        62008 => X"B8",  -- 184
        62009 => X"C2",  -- 194
        62010 => X"C4",  -- 196
        62011 => X"C7",  -- 199
        62012 => X"D2",  -- 210
        62013 => X"D7",  -- 215
        62014 => X"D5",  -- 213
        62015 => X"D6",  -- 214
        62016 => X"D5",  -- 213
        62017 => X"C3",  -- 195
        62018 => X"E0",  -- 224
        62019 => X"E1",  -- 225
        62020 => X"AD",  -- 173
        62021 => X"9C",  -- 156
        62022 => X"B7",  -- 183
        62023 => X"CF",  -- 207
        62024 => X"C8",  -- 200
        62025 => X"CF",  -- 207
        62026 => X"D8",  -- 216
        62027 => X"DC",  -- 220
        62028 => X"DC",  -- 220
        62029 => X"DA",  -- 218
        62030 => X"DB",  -- 219
        62031 => X"DC",  -- 220
        62032 => X"DB",  -- 219
        62033 => X"D2",  -- 210
        62034 => X"D0",  -- 208
        62035 => X"D1",  -- 209
        62036 => X"CE",  -- 206
        62037 => X"90",  -- 144
        62038 => X"40",  -- 64
        62039 => X"3D",  -- 61
        62040 => X"33",  -- 51
        62041 => X"2D",  -- 45
        62042 => X"2B",  -- 43
        62043 => X"2B",  -- 43
        62044 => X"2C",  -- 44
        62045 => X"28",  -- 40
        62046 => X"27",  -- 39
        62047 => X"28",  -- 40
        62048 => X"2C",  -- 44
        62049 => X"2D",  -- 45
        62050 => X"2D",  -- 45
        62051 => X"2D",  -- 45
        62052 => X"2C",  -- 44
        62053 => X"2A",  -- 42
        62054 => X"2A",  -- 42
        62055 => X"2A",  -- 42
        62056 => X"30",  -- 48
        62057 => X"34",  -- 52
        62058 => X"38",  -- 56
        62059 => X"3B",  -- 59
        62060 => X"3F",  -- 63
        62061 => X"48",  -- 72
        62062 => X"54",  -- 84
        62063 => X"5D",  -- 93
        62064 => X"5B",  -- 91
        62065 => X"63",  -- 99
        62066 => X"68",  -- 104
        62067 => X"5D",  -- 93
        62068 => X"5A",  -- 90
        62069 => X"6F",  -- 111
        62070 => X"85",  -- 133
        62071 => X"83",  -- 131
        62072 => X"85",  -- 133
        62073 => X"85",  -- 133
        62074 => X"6E",  -- 110
        62075 => X"63",  -- 99
        62076 => X"75",  -- 117
        62077 => X"75",  -- 117
        62078 => X"71",  -- 113
        62079 => X"7C",  -- 124
        62080 => X"53",  -- 83
        62081 => X"54",  -- 84
        62082 => X"55",  -- 85
        62083 => X"56",  -- 86
        62084 => X"58",  -- 88
        62085 => X"5B",  -- 91
        62086 => X"5F",  -- 95
        62087 => X"63",  -- 99
        62088 => X"60",  -- 96
        62089 => X"57",  -- 87
        62090 => X"4C",  -- 76
        62091 => X"4A",  -- 74
        62092 => X"53",  -- 83
        62093 => X"5B",  -- 91
        62094 => X"58",  -- 88
        62095 => X"50",  -- 80
        62096 => X"56",  -- 86
        62097 => X"67",  -- 103
        62098 => X"80",  -- 128
        62099 => X"74",  -- 116
        62100 => X"50",  -- 80
        62101 => X"4D",  -- 77
        62102 => X"54",  -- 84
        62103 => X"41",  -- 65
        62104 => X"3F",  -- 63
        62105 => X"55",  -- 85
        62106 => X"3D",  -- 61
        62107 => X"63",  -- 99
        62108 => X"9A",  -- 154
        62109 => X"8E",  -- 142
        62110 => X"79",  -- 121
        62111 => X"5E",  -- 94
        62112 => X"5B",  -- 91
        62113 => X"59",  -- 89
        62114 => X"90",  -- 144
        62115 => X"80",  -- 128
        62116 => X"79",  -- 121
        62117 => X"59",  -- 89
        62118 => X"66",  -- 102
        62119 => X"5C",  -- 92
        62120 => X"5B",  -- 91
        62121 => X"56",  -- 86
        62122 => X"5C",  -- 92
        62123 => X"6F",  -- 111
        62124 => X"66",  -- 102
        62125 => X"5B",  -- 91
        62126 => X"98",  -- 152
        62127 => X"8A",  -- 138
        62128 => X"5E",  -- 94
        62129 => X"52",  -- 82
        62130 => X"7A",  -- 122
        62131 => X"67",  -- 103
        62132 => X"5B",  -- 91
        62133 => X"85",  -- 133
        62134 => X"95",  -- 149
        62135 => X"72",  -- 114
        62136 => X"5C",  -- 92
        62137 => X"6B",  -- 107
        62138 => X"96",  -- 150
        62139 => X"4E",  -- 78
        62140 => X"6C",  -- 108
        62141 => X"7A",  -- 122
        62142 => X"6E",  -- 110
        62143 => X"79",  -- 121
        62144 => X"6E",  -- 110
        62145 => X"58",  -- 88
        62146 => X"49",  -- 73
        62147 => X"48",  -- 72
        62148 => X"67",  -- 103
        62149 => X"4A",  -- 74
        62150 => X"5D",  -- 93
        62151 => X"2A",  -- 42
        62152 => X"12",  -- 18
        62153 => X"14",  -- 20
        62154 => X"35",  -- 53
        62155 => X"1C",  -- 28
        62156 => X"1E",  -- 30
        62157 => X"1E",  -- 30
        62158 => X"23",  -- 35
        62159 => X"2B",  -- 43
        62160 => X"2E",  -- 46
        62161 => X"33",  -- 51
        62162 => X"37",  -- 55
        62163 => X"24",  -- 36
        62164 => X"20",  -- 32
        62165 => X"2D",  -- 45
        62166 => X"27",  -- 39
        62167 => X"23",  -- 35
        62168 => X"30",  -- 48
        62169 => X"2F",  -- 47
        62170 => X"34",  -- 52
        62171 => X"51",  -- 81
        62172 => X"6F",  -- 111
        62173 => X"5F",  -- 95
        62174 => X"38",  -- 56
        62175 => X"28",  -- 40
        62176 => X"2E",  -- 46
        62177 => X"30",  -- 48
        62178 => X"27",  -- 39
        62179 => X"29",  -- 41
        62180 => X"13",  -- 19
        62181 => X"1E",  -- 30
        62182 => X"42",  -- 66
        62183 => X"32",  -- 50
        62184 => X"15",  -- 21
        62185 => X"43",  -- 67
        62186 => X"4D",  -- 77
        62187 => X"4C",  -- 76
        62188 => X"49",  -- 73
        62189 => X"3F",  -- 63
        62190 => X"35",  -- 53
        62191 => X"2F",  -- 47
        62192 => X"27",  -- 39
        62193 => X"18",  -- 24
        62194 => X"57",  -- 87
        62195 => X"3B",  -- 59
        62196 => X"0D",  -- 13
        62197 => X"12",  -- 18
        62198 => X"67",  -- 103
        62199 => X"38",  -- 56
        62200 => X"4F",  -- 79
        62201 => X"66",  -- 102
        62202 => X"49",  -- 73
        62203 => X"58",  -- 88
        62204 => X"47",  -- 71
        62205 => X"5C",  -- 92
        62206 => X"84",  -- 132
        62207 => X"6F",  -- 111
        62208 => X"60",  -- 96
        62209 => X"84",  -- 132
        62210 => X"62",  -- 98
        62211 => X"8E",  -- 142
        62212 => X"88",  -- 136
        62213 => X"75",  -- 117
        62214 => X"85",  -- 133
        62215 => X"89",  -- 137
        62216 => X"51",  -- 81
        62217 => X"3B",  -- 59
        62218 => X"44",  -- 68
        62219 => X"4F",  -- 79
        62220 => X"39",  -- 57
        62221 => X"65",  -- 101
        62222 => X"B9",  -- 185
        62223 => X"6F",  -- 111
        62224 => X"36",  -- 54
        62225 => X"4A",  -- 74
        62226 => X"42",  -- 66
        62227 => X"48",  -- 72
        62228 => X"3D",  -- 61
        62229 => X"8B",  -- 139
        62230 => X"79",  -- 121
        62231 => X"7C",  -- 124
        62232 => X"50",  -- 80
        62233 => X"6E",  -- 110
        62234 => X"7A",  -- 122
        62235 => X"55",  -- 85
        62236 => X"62",  -- 98
        62237 => X"52",  -- 82
        62238 => X"2E",  -- 46
        62239 => X"4A",  -- 74
        62240 => X"43",  -- 67
        62241 => X"36",  -- 54
        62242 => X"28",  -- 40
        62243 => X"1B",  -- 27
        62244 => X"12",  -- 18
        62245 => X"0D",  -- 13
        62246 => X"11",  -- 17
        62247 => X"16",  -- 22
        62248 => X"16",  -- 22
        62249 => X"0C",  -- 12
        62250 => X"5B",  -- 91
        62251 => X"66",  -- 102
        62252 => X"13",  -- 19
        62253 => X"24",  -- 36
        62254 => X"0E",  -- 14
        62255 => X"15",  -- 21
        62256 => X"10",  -- 16
        62257 => X"17",  -- 23
        62258 => X"1D",  -- 29
        62259 => X"23",  -- 35
        62260 => X"2D",  -- 45
        62261 => X"3B",  -- 59
        62262 => X"43",  -- 67
        62263 => X"43",  -- 67
        62264 => X"3E",  -- 62
        62265 => X"3B",  -- 59
        62266 => X"3B",  -- 59
        62267 => X"37",  -- 55
        62268 => X"33",  -- 51
        62269 => X"32",  -- 50
        62270 => X"36",  -- 54
        62271 => X"3D",  -- 61
        62272 => X"44",  -- 68
        62273 => X"50",  -- 80
        62274 => X"61",  -- 97
        62275 => X"6B",  -- 107
        62276 => X"64",  -- 100
        62277 => X"54",  -- 84
        62278 => X"42",  -- 66
        62279 => X"37",  -- 55
        62280 => X"46",  -- 70
        62281 => X"48",  -- 72
        62282 => X"46",  -- 70
        62283 => X"3A",  -- 58
        62284 => X"30",  -- 48
        62285 => X"2D",  -- 45
        62286 => X"32",  -- 50
        62287 => X"36",  -- 54
        62288 => X"3D",  -- 61
        62289 => X"37",  -- 55
        62290 => X"81",  -- 129
        62291 => X"97",  -- 151
        62292 => X"96",  -- 150
        62293 => X"9F",  -- 159
        62294 => X"94",  -- 148
        62295 => X"92",  -- 146
        62296 => X"8D",  -- 141
        62297 => X"77",  -- 119
        62298 => X"8A",  -- 138
        62299 => X"7E",  -- 126
        62300 => X"68",  -- 104
        62301 => X"85",  -- 133
        62302 => X"85",  -- 133
        62303 => X"50",  -- 80
        62304 => X"0B",  -- 11
        62305 => X"12",  -- 18
        62306 => X"60",  -- 96
        62307 => X"87",  -- 135
        62308 => X"A0",  -- 160
        62309 => X"96",  -- 150
        62310 => X"A9",  -- 169
        62311 => X"AE",  -- 174
        62312 => X"9B",  -- 155
        62313 => X"A2",  -- 162
        62314 => X"A4",  -- 164
        62315 => X"AE",  -- 174
        62316 => X"70",  -- 112
        62317 => X"09",  -- 9
        62318 => X"00",  -- 0
        62319 => X"18",  -- 24
        62320 => X"5D",  -- 93
        62321 => X"9F",  -- 159
        62322 => X"A2",  -- 162
        62323 => X"60",  -- 96
        62324 => X"61",  -- 97
        62325 => X"B6",  -- 182
        62326 => X"AB",  -- 171
        62327 => X"AD",  -- 173
        62328 => X"BC",  -- 188
        62329 => X"C4",  -- 196
        62330 => X"C5",  -- 197
        62331 => X"C5",  -- 197
        62332 => X"CF",  -- 207
        62333 => X"D4",  -- 212
        62334 => X"D1",  -- 209
        62335 => X"D4",  -- 212
        62336 => X"D0",  -- 208
        62337 => X"CB",  -- 203
        62338 => X"D6",  -- 214
        62339 => X"E5",  -- 229
        62340 => X"C6",  -- 198
        62341 => X"A4",  -- 164
        62342 => X"B2",  -- 178
        62343 => X"C5",  -- 197
        62344 => X"C4",  -- 196
        62345 => X"CE",  -- 206
        62346 => X"D7",  -- 215
        62347 => X"DA",  -- 218
        62348 => X"DC",  -- 220
        62349 => X"E0",  -- 224
        62350 => X"E0",  -- 224
        62351 => X"DD",  -- 221
        62352 => X"DF",  -- 223
        62353 => X"D6",  -- 214
        62354 => X"D0",  -- 208
        62355 => X"D3",  -- 211
        62356 => X"CD",  -- 205
        62357 => X"8F",  -- 143
        62358 => X"45",  -- 69
        62359 => X"40",  -- 64
        62360 => X"33",  -- 51
        62361 => X"2E",  -- 46
        62362 => X"2D",  -- 45
        62363 => X"2E",  -- 46
        62364 => X"31",  -- 49
        62365 => X"2D",  -- 45
        62366 => X"29",  -- 41
        62367 => X"29",  -- 41
        62368 => X"2F",  -- 47
        62369 => X"2F",  -- 47
        62370 => X"30",  -- 48
        62371 => X"2E",  -- 46
        62372 => X"2C",  -- 44
        62373 => X"2C",  -- 44
        62374 => X"30",  -- 48
        62375 => X"33",  -- 51
        62376 => X"33",  -- 51
        62377 => X"37",  -- 55
        62378 => X"3C",  -- 60
        62379 => X"3F",  -- 63
        62380 => X"42",  -- 66
        62381 => X"49",  -- 73
        62382 => X"55",  -- 85
        62383 => X"5F",  -- 95
        62384 => X"5B",  -- 91
        62385 => X"5D",  -- 93
        62386 => X"5C",  -- 92
        62387 => X"54",  -- 84
        62388 => X"55",  -- 85
        62389 => X"6E",  -- 110
        62390 => X"84",  -- 132
        62391 => X"84",  -- 132
        62392 => X"84",  -- 132
        62393 => X"76",  -- 118
        62394 => X"5C",  -- 92
        62395 => X"5C",  -- 92
        62396 => X"70",  -- 112
        62397 => X"74",  -- 116
        62398 => X"6C",  -- 108
        62399 => X"75",  -- 117
        62400 => X"5F",  -- 95
        62401 => X"61",  -- 97
        62402 => X"63",  -- 99
        62403 => X"65",  -- 101
        62404 => X"68",  -- 104
        62405 => X"6B",  -- 107
        62406 => X"6F",  -- 111
        62407 => X"72",  -- 114
        62408 => X"7C",  -- 124
        62409 => X"6F",  -- 111
        62410 => X"5F",  -- 95
        62411 => X"58",  -- 88
        62412 => X"5C",  -- 92
        62413 => X"64",  -- 100
        62414 => X"68",  -- 104
        62415 => X"68",  -- 104
        62416 => X"74",  -- 116
        62417 => X"8E",  -- 142
        62418 => X"75",  -- 117
        62419 => X"4A",  -- 74
        62420 => X"48",  -- 72
        62421 => X"4D",  -- 77
        62422 => X"4A",  -- 74
        62423 => X"55",  -- 85
        62424 => X"56",  -- 86
        62425 => X"4E",  -- 78
        62426 => X"51",  -- 81
        62427 => X"9B",  -- 155
        62428 => X"95",  -- 149
        62429 => X"57",  -- 87
        62430 => X"64",  -- 100
        62431 => X"5F",  -- 95
        62432 => X"66",  -- 102
        62433 => X"81",  -- 129
        62434 => X"93",  -- 147
        62435 => X"6D",  -- 109
        62436 => X"60",  -- 96
        62437 => X"69",  -- 105
        62438 => X"59",  -- 89
        62439 => X"59",  -- 89
        62440 => X"58",  -- 88
        62441 => X"53",  -- 83
        62442 => X"70",  -- 112
        62443 => X"6F",  -- 111
        62444 => X"54",  -- 84
        62445 => X"91",  -- 145
        62446 => X"9E",  -- 158
        62447 => X"53",  -- 83
        62448 => X"4D",  -- 77
        62449 => X"72",  -- 114
        62450 => X"72",  -- 114
        62451 => X"44",  -- 68
        62452 => X"6B",  -- 107
        62453 => X"8D",  -- 141
        62454 => X"6A",  -- 106
        62455 => X"6D",  -- 109
        62456 => X"6E",  -- 110
        62457 => X"7D",  -- 125
        62458 => X"77",  -- 119
        62459 => X"4A",  -- 74
        62460 => X"86",  -- 134
        62461 => X"78",  -- 120
        62462 => X"7E",  -- 126
        62463 => X"64",  -- 100
        62464 => X"4F",  -- 79
        62465 => X"4F",  -- 79
        62466 => X"42",  -- 66
        62467 => X"6C",  -- 108
        62468 => X"54",  -- 84
        62469 => X"4F",  -- 79
        62470 => X"5D",  -- 93
        62471 => X"22",  -- 34
        62472 => X"24",  -- 36
        62473 => X"2C",  -- 44
        62474 => X"49",  -- 73
        62475 => X"29",  -- 41
        62476 => X"38",  -- 56
        62477 => X"32",  -- 50
        62478 => X"3C",  -- 60
        62479 => X"41",  -- 65
        62480 => X"44",  -- 68
        62481 => X"3D",  -- 61
        62482 => X"3E",  -- 62
        62483 => X"36",  -- 54
        62484 => X"37",  -- 55
        62485 => X"3D",  -- 61
        62486 => X"31",  -- 49
        62487 => X"2F",  -- 47
        62488 => X"3D",  -- 61
        62489 => X"3C",  -- 60
        62490 => X"40",  -- 64
        62491 => X"5B",  -- 91
        62492 => X"6A",  -- 106
        62493 => X"48",  -- 72
        62494 => X"34",  -- 52
        62495 => X"51",  -- 81
        62496 => X"38",  -- 56
        62497 => X"36",  -- 54
        62498 => X"28",  -- 40
        62499 => X"36",  -- 54
        62500 => X"1E",  -- 30
        62501 => X"22",  -- 34
        62502 => X"3C",  -- 60
        62503 => X"31",  -- 49
        62504 => X"1A",  -- 26
        62505 => X"47",  -- 71
        62506 => X"41",  -- 65
        62507 => X"5E",  -- 94
        62508 => X"3F",  -- 63
        62509 => X"44",  -- 68
        62510 => X"22",  -- 34
        62511 => X"33",  -- 51
        62512 => X"33",  -- 51
        62513 => X"36",  -- 54
        62514 => X"37",  -- 55
        62515 => X"43",  -- 67
        62516 => X"38",  -- 56
        62517 => X"10",  -- 16
        62518 => X"3B",  -- 59
        62519 => X"69",  -- 105
        62520 => X"45",  -- 69
        62521 => X"5B",  -- 91
        62522 => X"65",  -- 101
        62523 => X"3E",  -- 62
        62524 => X"61",  -- 97
        62525 => X"65",  -- 101
        62526 => X"56",  -- 86
        62527 => X"7E",  -- 126
        62528 => X"58",  -- 88
        62529 => X"69",  -- 105
        62530 => X"7B",  -- 123
        62531 => X"68",  -- 104
        62532 => X"96",  -- 150
        62533 => X"88",  -- 136
        62534 => X"39",  -- 57
        62535 => X"7B",  -- 123
        62536 => X"B6",  -- 182
        62537 => X"6A",  -- 106
        62538 => X"3A",  -- 58
        62539 => X"44",  -- 68
        62540 => X"37",  -- 55
        62541 => X"3C",  -- 60
        62542 => X"8D",  -- 141
        62543 => X"AA",  -- 170
        62544 => X"61",  -- 97
        62545 => X"34",  -- 52
        62546 => X"50",  -- 80
        62547 => X"45",  -- 69
        62548 => X"51",  -- 81
        62549 => X"3C",  -- 60
        62550 => X"82",  -- 130
        62551 => X"86",  -- 134
        62552 => X"81",  -- 129
        62553 => X"46",  -- 70
        62554 => X"79",  -- 121
        62555 => X"75",  -- 117
        62556 => X"56",  -- 86
        62557 => X"55",  -- 85
        62558 => X"41",  -- 65
        62559 => X"45",  -- 69
        62560 => X"3B",  -- 59
        62561 => X"26",  -- 38
        62562 => X"14",  -- 20
        62563 => X"10",  -- 16
        62564 => X"0F",  -- 15
        62565 => X"0A",  -- 10
        62566 => X"0C",  -- 12
        62567 => X"14",  -- 20
        62568 => X"16",  -- 22
        62569 => X"0A",  -- 10
        62570 => X"1B",  -- 27
        62571 => X"42",  -- 66
        62572 => X"69",  -- 105
        62573 => X"1C",  -- 28
        62574 => X"0D",  -- 13
        62575 => X"10",  -- 16
        62576 => X"1D",  -- 29
        62577 => X"25",  -- 37
        62578 => X"2B",  -- 43
        62579 => X"2E",  -- 46
        62580 => X"33",  -- 51
        62581 => X"39",  -- 57
        62582 => X"3B",  -- 59
        62583 => X"3A",  -- 58
        62584 => X"39",  -- 57
        62585 => X"3A",  -- 58
        62586 => X"39",  -- 57
        62587 => X"36",  -- 54
        62588 => X"33",  -- 51
        62589 => X"35",  -- 53
        62590 => X"3A",  -- 58
        62591 => X"40",  -- 64
        62592 => X"3E",  -- 62
        62593 => X"4A",  -- 74
        62594 => X"5D",  -- 93
        62595 => X"69",  -- 105
        62596 => X"66",  -- 102
        62597 => X"55",  -- 85
        62598 => X"44",  -- 68
        62599 => X"3C",  -- 60
        62600 => X"4E",  -- 78
        62601 => X"51",  -- 81
        62602 => X"4D",  -- 77
        62603 => X"40",  -- 64
        62604 => X"35",  -- 53
        62605 => X"32",  -- 50
        62606 => X"35",  -- 53
        62607 => X"38",  -- 56
        62608 => X"31",  -- 49
        62609 => X"5B",  -- 91
        62610 => X"9C",  -- 156
        62611 => X"87",  -- 135
        62612 => X"91",  -- 145
        62613 => X"A1",  -- 161
        62614 => X"96",  -- 150
        62615 => X"8A",  -- 138
        62616 => X"7F",  -- 127
        62617 => X"72",  -- 114
        62618 => X"8F",  -- 143
        62619 => X"8F",  -- 143
        62620 => X"7B",  -- 123
        62621 => X"83",  -- 131
        62622 => X"64",  -- 100
        62623 => X"21",  -- 33
        62624 => X"07",  -- 7
        62625 => X"38",  -- 56
        62626 => X"95",  -- 149
        62627 => X"89",  -- 137
        62628 => X"A8",  -- 168
        62629 => X"98",  -- 152
        62630 => X"BB",  -- 187
        62631 => X"AF",  -- 175
        62632 => X"AA",  -- 170
        62633 => X"A9",  -- 169
        62634 => X"A1",  -- 161
        62635 => X"A0",  -- 160
        62636 => X"37",  -- 55
        62637 => X"01",  -- 1
        62638 => X"00",  -- 0
        62639 => X"26",  -- 38
        62640 => X"6B",  -- 107
        62641 => X"A0",  -- 160
        62642 => X"9C",  -- 156
        62643 => X"50",  -- 80
        62644 => X"37",  -- 55
        62645 => X"A8",  -- 168
        62646 => X"B5",  -- 181
        62647 => X"BA",  -- 186
        62648 => X"BD",  -- 189
        62649 => X"C3",  -- 195
        62650 => X"C2",  -- 194
        62651 => X"C2",  -- 194
        62652 => X"CC",  -- 204
        62653 => X"CF",  -- 207
        62654 => X"CA",  -- 202
        62655 => X"CB",  -- 203
        62656 => X"D0",  -- 208
        62657 => X"D6",  -- 214
        62658 => X"C6",  -- 198
        62659 => X"D2",  -- 210
        62660 => X"D3",  -- 211
        62661 => X"B9",  -- 185
        62662 => X"B5",  -- 181
        62663 => X"B0",  -- 176
        62664 => X"C7",  -- 199
        62665 => X"C8",  -- 200
        62666 => X"CC",  -- 204
        62667 => X"D2",  -- 210
        62668 => X"D8",  -- 216
        62669 => X"DC",  -- 220
        62670 => X"DE",  -- 222
        62671 => X"DD",  -- 221
        62672 => X"DF",  -- 223
        62673 => X"D6",  -- 214
        62674 => X"D1",  -- 209
        62675 => X"D5",  -- 213
        62676 => X"CB",  -- 203
        62677 => X"8B",  -- 139
        62678 => X"4B",  -- 75
        62679 => X"41",  -- 65
        62680 => X"35",  -- 53
        62681 => X"31",  -- 49
        62682 => X"30",  -- 48
        62683 => X"34",  -- 52
        62684 => X"37",  -- 55
        62685 => X"35",  -- 53
        62686 => X"31",  -- 49
        62687 => X"31",  -- 49
        62688 => X"2E",  -- 46
        62689 => X"31",  -- 49
        62690 => X"32",  -- 50
        62691 => X"31",  -- 49
        62692 => X"2C",  -- 44
        62693 => X"2B",  -- 43
        62694 => X"2F",  -- 47
        62695 => X"35",  -- 53
        62696 => X"34",  -- 52
        62697 => X"39",  -- 57
        62698 => X"3F",  -- 63
        62699 => X"41",  -- 65
        62700 => X"44",  -- 68
        62701 => X"49",  -- 73
        62702 => X"52",  -- 82
        62703 => X"59",  -- 89
        62704 => X"55",  -- 85
        62705 => X"53",  -- 83
        62706 => X"52",  -- 82
        62707 => X"4F",  -- 79
        62708 => X"53",  -- 83
        62709 => X"6B",  -- 107
        62710 => X"80",  -- 128
        62711 => X"7E",  -- 126
        62712 => X"7C",  -- 124
        62713 => X"67",  -- 103
        62714 => X"51",  -- 81
        62715 => X"56",  -- 86
        62716 => X"6B",  -- 107
        62717 => X"6C",  -- 108
        62718 => X"66",  -- 102
        62719 => X"6C",  -- 108
        62720 => X"71",  -- 113
        62721 => X"74",  -- 116
        62722 => X"77",  -- 119
        62723 => X"79",  -- 121
        62724 => X"7A",  -- 122
        62725 => X"7B",  -- 123
        62726 => X"7D",  -- 125
        62727 => X"7E",  -- 126
        62728 => X"7B",  -- 123
        62729 => X"78",  -- 120
        62730 => X"76",  -- 118
        62731 => X"75",  -- 117
        62732 => X"77",  -- 119
        62733 => X"7A",  -- 122
        62734 => X"7D",  -- 125
        62735 => X"7F",  -- 127
        62736 => X"96",  -- 150
        62737 => X"70",  -- 112
        62738 => X"67",  -- 103
        62739 => X"68",  -- 104
        62740 => X"59",  -- 89
        62741 => X"5D",  -- 93
        62742 => X"68",  -- 104
        62743 => X"5D",  -- 93
        62744 => X"59",  -- 89
        62745 => X"68",  -- 104
        62746 => X"93",  -- 147
        62747 => X"64",  -- 100
        62748 => X"46",  -- 70
        62749 => X"68",  -- 104
        62750 => X"5C",  -- 92
        62751 => X"5C",  -- 92
        62752 => X"76",  -- 118
        62753 => X"90",  -- 144
        62754 => X"52",  -- 82
        62755 => X"83",  -- 131
        62756 => X"51",  -- 81
        62757 => X"5E",  -- 94
        62758 => X"55",  -- 85
        62759 => X"5E",  -- 94
        62760 => X"5B",  -- 91
        62761 => X"4A",  -- 74
        62762 => X"84",  -- 132
        62763 => X"55",  -- 85
        62764 => X"69",  -- 105
        62765 => X"A9",  -- 169
        62766 => X"64",  -- 100
        62767 => X"46",  -- 70
        62768 => X"62",  -- 98
        62769 => X"7B",  -- 123
        62770 => X"46",  -- 70
        62771 => X"65",  -- 101
        62772 => X"8C",  -- 140
        62773 => X"6A",  -- 106
        62774 => X"6A",  -- 106
        62775 => X"6F",  -- 111
        62776 => X"65",  -- 101
        62777 => X"7F",  -- 127
        62778 => X"57",  -- 87
        62779 => X"70",  -- 112
        62780 => X"74",  -- 116
        62781 => X"76",  -- 118
        62782 => X"73",  -- 115
        62783 => X"61",  -- 97
        62784 => X"3E",  -- 62
        62785 => X"3E",  -- 62
        62786 => X"63",  -- 99
        62787 => X"5E",  -- 94
        62788 => X"51",  -- 81
        62789 => X"69",  -- 105
        62790 => X"3D",  -- 61
        62791 => X"3E",  -- 62
        62792 => X"36",  -- 54
        62793 => X"3B",  -- 59
        62794 => X"52",  -- 82
        62795 => X"3C",  -- 60
        62796 => X"50",  -- 80
        62797 => X"45",  -- 69
        62798 => X"55",  -- 85
        62799 => X"5B",  -- 91
        62800 => X"56",  -- 86
        62801 => X"3A",  -- 58
        62802 => X"3A",  -- 58
        62803 => X"4C",  -- 76
        62804 => X"5C",  -- 92
        62805 => X"56",  -- 86
        62806 => X"3E",  -- 62
        62807 => X"3C",  -- 60
        62808 => X"4D",  -- 77
        62809 => X"50",  -- 80
        62810 => X"4B",  -- 75
        62811 => X"50",  -- 80
        62812 => X"52",  -- 82
        62813 => X"39",  -- 57
        62814 => X"37",  -- 55
        62815 => X"5D",  -- 93
        62816 => X"40",  -- 64
        62817 => X"46",  -- 70
        62818 => X"38",  -- 56
        62819 => X"4D",  -- 77
        62820 => X"31",  -- 49
        62821 => X"27",  -- 39
        62822 => X"3C",  -- 60
        62823 => X"4A",  -- 74
        62824 => X"53",  -- 83
        62825 => X"67",  -- 103
        62826 => X"51",  -- 81
        62827 => X"66",  -- 102
        62828 => X"50",  -- 80
        62829 => X"64",  -- 100
        62830 => X"32",  -- 50
        62831 => X"2D",  -- 45
        62832 => X"3F",  -- 63
        62833 => X"58",  -- 88
        62834 => X"44",  -- 68
        62835 => X"5A",  -- 90
        62836 => X"53",  -- 83
        62837 => X"2D",  -- 45
        62838 => X"32",  -- 50
        62839 => X"63",  -- 99
        62840 => X"56",  -- 86
        62841 => X"3D",  -- 61
        62842 => X"73",  -- 115
        62843 => X"59",  -- 89
        62844 => X"5A",  -- 90
        62845 => X"5C",  -- 92
        62846 => X"47",  -- 71
        62847 => X"67",  -- 103
        62848 => X"6F",  -- 111
        62849 => X"5B",  -- 91
        62850 => X"59",  -- 89
        62851 => X"6F",  -- 111
        62852 => X"63",  -- 99
        62853 => X"A7",  -- 167
        62854 => X"48",  -- 72
        62855 => X"40",  -- 64
        62856 => X"67",  -- 103
        62857 => X"9C",  -- 156
        62858 => X"63",  -- 99
        62859 => X"4A",  -- 74
        62860 => X"46",  -- 70
        62861 => X"39",  -- 57
        62862 => X"67",  -- 103
        62863 => X"53",  -- 83
        62864 => X"8C",  -- 140
        62865 => X"4F",  -- 79
        62866 => X"43",  -- 67
        62867 => X"58",  -- 88
        62868 => X"48",  -- 72
        62869 => X"59",  -- 89
        62870 => X"45",  -- 69
        62871 => X"74",  -- 116
        62872 => X"7C",  -- 124
        62873 => X"90",  -- 144
        62874 => X"37",  -- 55
        62875 => X"85",  -- 133
        62876 => X"6E",  -- 110
        62877 => X"50",  -- 80
        62878 => X"4D",  -- 77
        62879 => X"3F",  -- 63
        62880 => X"2D",  -- 45
        62881 => X"18",  -- 24
        62882 => X"0B",  -- 11
        62883 => X"0D",  -- 13
        62884 => X"0F",  -- 15
        62885 => X"0B",  -- 11
        62886 => X"0D",  -- 13
        62887 => X"14",  -- 20
        62888 => X"11",  -- 17
        62889 => X"19",  -- 25
        62890 => X"09",  -- 9
        62891 => X"17",  -- 23
        62892 => X"2A",  -- 42
        62893 => X"4F",  -- 79
        62894 => X"1B",  -- 27
        62895 => X"14",  -- 20
        62896 => X"1C",  -- 28
        62897 => X"21",  -- 33
        62898 => X"25",  -- 37
        62899 => X"24",  -- 36
        62900 => X"24",  -- 36
        62901 => X"23",  -- 35
        62902 => X"22",  -- 34
        62903 => X"21",  -- 33
        62904 => X"1D",  -- 29
        62905 => X"1C",  -- 28
        62906 => X"1C",  -- 28
        62907 => X"1D",  -- 29
        62908 => X"21",  -- 33
        62909 => X"28",  -- 40
        62910 => X"2E",  -- 46
        62911 => X"31",  -- 49
        62912 => X"34",  -- 52
        62913 => X"40",  -- 64
        62914 => X"53",  -- 83
        62915 => X"63",  -- 99
        62916 => X"62",  -- 98
        62917 => X"54",  -- 84
        62918 => X"46",  -- 70
        62919 => X"41",  -- 65
        62920 => X"52",  -- 82
        62921 => X"52",  -- 82
        62922 => X"4C",  -- 76
        62923 => X"3F",  -- 63
        62924 => X"34",  -- 52
        62925 => X"33",  -- 51
        62926 => X"35",  -- 53
        62927 => X"39",  -- 57
        62928 => X"39",  -- 57
        62929 => X"84",  -- 132
        62930 => X"8C",  -- 140
        62931 => X"6E",  -- 110
        62932 => X"95",  -- 149
        62933 => X"9A",  -- 154
        62934 => X"8D",  -- 141
        62935 => X"7A",  -- 122
        62936 => X"78",  -- 120
        62937 => X"76",  -- 118
        62938 => X"87",  -- 135
        62939 => X"8D",  -- 141
        62940 => X"89",  -- 137
        62941 => X"74",  -- 116
        62942 => X"38",  -- 56
        62943 => X"06",  -- 6
        62944 => X"0C",  -- 12
        62945 => X"56",  -- 86
        62946 => X"95",  -- 149
        62947 => X"A3",  -- 163
        62948 => X"A5",  -- 165
        62949 => X"A3",  -- 163
        62950 => X"B1",  -- 177
        62951 => X"BA",  -- 186
        62952 => X"B1",  -- 177
        62953 => X"9C",  -- 156
        62954 => X"9B",  -- 155
        62955 => X"74",  -- 116
        62956 => X"0A",  -- 10
        62957 => X"03",  -- 3
        62958 => X"00",  -- 0
        62959 => X"26",  -- 38
        62960 => X"6D",  -- 109
        62961 => X"93",  -- 147
        62962 => X"9B",  -- 155
        62963 => X"58",  -- 88
        62964 => X"20",  -- 32
        62965 => X"8F",  -- 143
        62966 => X"BF",  -- 191
        62967 => X"C4",  -- 196
        62968 => X"B8",  -- 184
        62969 => X"BF",  -- 191
        62970 => X"BD",  -- 189
        62971 => X"BC",  -- 188
        62972 => X"C6",  -- 198
        62973 => X"CA",  -- 202
        62974 => X"C5",  -- 197
        62975 => X"C3",  -- 195
        62976 => X"D1",  -- 209
        62977 => X"D5",  -- 213
        62978 => X"B8",  -- 184
        62979 => X"C2",  -- 194
        62980 => X"D3",  -- 211
        62981 => X"BC",  -- 188
        62982 => X"AE",  -- 174
        62983 => X"A6",  -- 166
        62984 => X"C5",  -- 197
        62985 => X"BE",  -- 190
        62986 => X"BF",  -- 191
        62987 => X"CA",  -- 202
        62988 => X"D3",  -- 211
        62989 => X"D2",  -- 210
        62990 => X"D0",  -- 208
        62991 => X"D3",  -- 211
        62992 => X"D7",  -- 215
        62993 => X"D1",  -- 209
        62994 => X"CD",  -- 205
        62995 => X"D5",  -- 213
        62996 => X"C1",  -- 193
        62997 => X"7D",  -- 125
        62998 => X"4A",  -- 74
        62999 => X"40",  -- 64
        63000 => X"38",  -- 56
        63001 => X"33",  -- 51
        63002 => X"31",  -- 49
        63003 => X"38",  -- 56
        63004 => X"3C",  -- 60
        63005 => X"3D",  -- 61
        63006 => X"3C",  -- 60
        63007 => X"3B",  -- 59
        63008 => X"33",  -- 51
        63009 => X"3A",  -- 58
        63010 => X"3E",  -- 62
        63011 => X"3B",  -- 59
        63012 => X"34",  -- 52
        63013 => X"2F",  -- 47
        63014 => X"32",  -- 50
        63015 => X"35",  -- 53
        63016 => X"37",  -- 55
        63017 => X"3B",  -- 59
        63018 => X"40",  -- 64
        63019 => X"42",  -- 66
        63020 => X"45",  -- 69
        63021 => X"47",  -- 71
        63022 => X"4B",  -- 75
        63023 => X"4F",  -- 79
        63024 => X"4C",  -- 76
        63025 => X"48",  -- 72
        63026 => X"49",  -- 73
        63027 => X"4B",  -- 75
        63028 => X"51",  -- 81
        63029 => X"63",  -- 99
        63030 => X"73",  -- 115
        63031 => X"70",  -- 112
        63032 => X"6B",  -- 107
        63033 => X"59",  -- 89
        63034 => X"4C",  -- 76
        63035 => X"54",  -- 84
        63036 => X"63",  -- 99
        63037 => X"63",  -- 99
        63038 => X"5F",  -- 95
        63039 => X"64",  -- 100
        63040 => X"76",  -- 118
        63041 => X"78",  -- 120
        63042 => X"7B",  -- 123
        63043 => X"7C",  -- 124
        63044 => X"7B",  -- 123
        63045 => X"7A",  -- 122
        63046 => X"79",  -- 121
        63047 => X"79",  -- 121
        63048 => X"76",  -- 118
        63049 => X"74",  -- 116
        63050 => X"73",  -- 115
        63051 => X"73",  -- 115
        63052 => X"72",  -- 114
        63053 => X"74",  -- 116
        63054 => X"7B",  -- 123
        63055 => X"83",  -- 131
        63056 => X"64",  -- 100
        63057 => X"74",  -- 116
        63058 => X"6D",  -- 109
        63059 => X"64",  -- 100
        63060 => X"6A",  -- 106
        63061 => X"61",  -- 97
        63062 => X"5D",  -- 93
        63063 => X"72",  -- 114
        63064 => X"6F",  -- 111
        63065 => X"70",  -- 112
        63066 => X"71",  -- 113
        63067 => X"56",  -- 86
        63068 => X"5C",  -- 92
        63069 => X"5E",  -- 94
        63070 => X"4B",  -- 75
        63071 => X"79",  -- 121
        63072 => X"80",  -- 128
        63073 => X"63",  -- 99
        63074 => X"62",  -- 98
        63075 => X"78",  -- 120
        63076 => X"51",  -- 81
        63077 => X"50",  -- 80
        63078 => X"5B",  -- 91
        63079 => X"55",  -- 85
        63080 => X"53",  -- 83
        63081 => X"65",  -- 101
        63082 => X"67",  -- 103
        63083 => X"56",  -- 86
        63084 => X"96",  -- 150
        63085 => X"67",  -- 103
        63086 => X"45",  -- 69
        63087 => X"5E",  -- 94
        63088 => X"74",  -- 116
        63089 => X"51",  -- 81
        63090 => X"57",  -- 87
        63091 => X"8A",  -- 138
        63092 => X"79",  -- 121
        63093 => X"70",  -- 112
        63094 => X"7D",  -- 125
        63095 => X"62",  -- 98
        63096 => X"71",  -- 113
        63097 => X"52",  -- 82
        63098 => X"6A",  -- 106
        63099 => X"85",  -- 133
        63100 => X"5B",  -- 91
        63101 => X"6C",  -- 108
        63102 => X"72",  -- 114
        63103 => X"3D",  -- 61
        63104 => X"45",  -- 69
        63105 => X"54",  -- 84
        63106 => X"66",  -- 102
        63107 => X"3A",  -- 58
        63108 => X"70",  -- 112
        63109 => X"58",  -- 88
        63110 => X"34",  -- 52
        63111 => X"4B",  -- 75
        63112 => X"46",  -- 70
        63113 => X"44",  -- 68
        63114 => X"51",  -- 81
        63115 => X"47",  -- 71
        63116 => X"52",  -- 82
        63117 => X"48",  -- 72
        63118 => X"56",  -- 86
        63119 => X"57",  -- 87
        63120 => X"4D",  -- 77
        63121 => X"3F",  -- 63
        63122 => X"4D",  -- 77
        63123 => X"5D",  -- 93
        63124 => X"60",  -- 96
        63125 => X"51",  -- 81
        63126 => X"42",  -- 66
        63127 => X"4D",  -- 77
        63128 => X"58",  -- 88
        63129 => X"5B",  -- 91
        63130 => X"4B",  -- 75
        63131 => X"3D",  -- 61
        63132 => X"41",  -- 65
        63133 => X"3F",  -- 63
        63134 => X"3B",  -- 59
        63135 => X"43",  -- 67
        63136 => X"4E",  -- 78
        63137 => X"57",  -- 87
        63138 => X"39",  -- 57
        63139 => X"57",  -- 87
        63140 => X"51",  -- 81
        63141 => X"4E",  -- 78
        63142 => X"52",  -- 82
        63143 => X"65",  -- 101
        63144 => X"5F",  -- 95
        63145 => X"6A",  -- 106
        63146 => X"71",  -- 113
        63147 => X"63",  -- 99
        63148 => X"64",  -- 100
        63149 => X"77",  -- 119
        63150 => X"64",  -- 100
        63151 => X"4D",  -- 77
        63152 => X"69",  -- 105
        63153 => X"53",  -- 83
        63154 => X"66",  -- 102
        63155 => X"78",  -- 120
        63156 => X"53",  -- 83
        63157 => X"39",  -- 57
        63158 => X"4F",  -- 79
        63159 => X"50",  -- 80
        63160 => X"59",  -- 89
        63161 => X"45",  -- 69
        63162 => X"58",  -- 88
        63163 => X"73",  -- 115
        63164 => X"52",  -- 82
        63165 => X"54",  -- 84
        63166 => X"4F",  -- 79
        63167 => X"56",  -- 86
        63168 => X"83",  -- 131
        63169 => X"59",  -- 89
        63170 => X"46",  -- 70
        63171 => X"5A",  -- 90
        63172 => X"70",  -- 112
        63173 => X"62",  -- 98
        63174 => X"91",  -- 145
        63175 => X"47",  -- 71
        63176 => X"47",  -- 71
        63177 => X"69",  -- 105
        63178 => X"AD",  -- 173
        63179 => X"63",  -- 99
        63180 => X"40",  -- 64
        63181 => X"4B",  -- 75
        63182 => X"45",  -- 69
        63183 => X"83",  -- 131
        63184 => X"69",  -- 105
        63185 => X"8E",  -- 142
        63186 => X"3C",  -- 60
        63187 => X"48",  -- 72
        63188 => X"5E",  -- 94
        63189 => X"48",  -- 72
        63190 => X"51",  -- 81
        63191 => X"4C",  -- 76
        63192 => X"86",  -- 134
        63193 => X"58",  -- 88
        63194 => X"83",  -- 131
        63195 => X"50",  -- 80
        63196 => X"7C",  -- 124
        63197 => X"69",  -- 105
        63198 => X"4F",  -- 79
        63199 => X"31",  -- 49
        63200 => X"1E",  -- 30
        63201 => X"12",  -- 18
        63202 => X"0A",  -- 10
        63203 => X"11",  -- 17
        63204 => X"16",  -- 22
        63205 => X"12",  -- 18
        63206 => X"11",  -- 17
        63207 => X"17",  -- 23
        63208 => X"1A",  -- 26
        63209 => X"12",  -- 18
        63210 => X"15",  -- 21
        63211 => X"1E",  -- 30
        63212 => X"14",  -- 20
        63213 => X"1A",  -- 26
        63214 => X"70",  -- 112
        63215 => X"36",  -- 54
        63216 => X"16",  -- 22
        63217 => X"18",  -- 24
        63218 => X"17",  -- 23
        63219 => X"16",  -- 22
        63220 => X"16",  -- 22
        63221 => X"15",  -- 21
        63222 => X"14",  -- 20
        63223 => X"11",  -- 17
        63224 => X"13",  -- 19
        63225 => X"13",  -- 19
        63226 => X"13",  -- 19
        63227 => X"16",  -- 22
        63228 => X"1F",  -- 31
        63229 => X"2A",  -- 42
        63230 => X"2E",  -- 46
        63231 => X"2C",  -- 44
        63232 => X"2C",  -- 44
        63233 => X"34",  -- 52
        63234 => X"47",  -- 71
        63235 => X"58",  -- 88
        63236 => X"5C",  -- 92
        63237 => X"54",  -- 84
        63238 => X"4E",  -- 78
        63239 => X"4F",  -- 79
        63240 => X"5C",  -- 92
        63241 => X"57",  -- 87
        63242 => X"49",  -- 73
        63243 => X"3B",  -- 59
        63244 => X"31",  -- 49
        63245 => X"31",  -- 49
        63246 => X"34",  -- 52
        63247 => X"35",  -- 53
        63248 => X"46",  -- 70
        63249 => X"81",  -- 129
        63250 => X"5D",  -- 93
        63251 => X"62",  -- 98
        63252 => X"9A",  -- 154
        63253 => X"8C",  -- 140
        63254 => X"83",  -- 131
        63255 => X"74",  -- 116
        63256 => X"76",  -- 118
        63257 => X"74",  -- 116
        63258 => X"74",  -- 116
        63259 => X"75",  -- 117
        63260 => X"7D",  -- 125
        63261 => X"5E",  -- 94
        63262 => X"21",  -- 33
        63263 => X"0E",  -- 14
        63264 => X"15",  -- 21
        63265 => X"6B",  -- 107
        63266 => X"9E",  -- 158
        63267 => X"99",  -- 153
        63268 => X"A6",  -- 166
        63269 => X"A3",  -- 163
        63270 => X"AC",  -- 172
        63271 => X"9F",  -- 159
        63272 => X"AB",  -- 171
        63273 => X"8C",  -- 140
        63274 => X"9E",  -- 158
        63275 => X"51",  -- 81
        63276 => X"02",  -- 2
        63277 => X"06",  -- 6
        63278 => X"07",  -- 7
        63279 => X"18",  -- 24
        63280 => X"6D",  -- 109
        63281 => X"8D",  -- 141
        63282 => X"97",  -- 151
        63283 => X"60",  -- 96
        63284 => X"16",  -- 22
        63285 => X"5F",  -- 95
        63286 => X"AC",  -- 172
        63287 => X"C2",  -- 194
        63288 => X"BA",  -- 186
        63289 => X"BE",  -- 190
        63290 => X"B9",  -- 185
        63291 => X"B8",  -- 184
        63292 => X"C3",  -- 195
        63293 => X"C8",  -- 200
        63294 => X"C4",  -- 196
        63295 => X"C4",  -- 196
        63296 => X"CE",  -- 206
        63297 => X"C8",  -- 200
        63298 => X"B2",  -- 178
        63299 => X"BF",  -- 191
        63300 => X"CF",  -- 207
        63301 => X"AF",  -- 175
        63302 => X"97",  -- 151
        63303 => X"9E",  -- 158
        63304 => X"BE",  -- 190
        63305 => X"BD",  -- 189
        63306 => X"C0",  -- 192
        63307 => X"C7",  -- 199
        63308 => X"CC",  -- 204
        63309 => X"CB",  -- 203
        63310 => X"C9",  -- 201
        63311 => X"CA",  -- 202
        63312 => X"CD",  -- 205
        63313 => X"CE",  -- 206
        63314 => X"C9",  -- 201
        63315 => X"CF",  -- 207
        63316 => X"AE",  -- 174
        63317 => X"67",  -- 103
        63318 => X"42",  -- 66
        63319 => X"3F",  -- 63
        63320 => X"3A",  -- 58
        63321 => X"33",  -- 51
        63322 => X"2F",  -- 47
        63323 => X"37",  -- 55
        63324 => X"3F",  -- 63
        63325 => X"42",  -- 66
        63326 => X"45",  -- 69
        63327 => X"46",  -- 70
        63328 => X"40",  -- 64
        63329 => X"48",  -- 72
        63330 => X"50",  -- 80
        63331 => X"4C",  -- 76
        63332 => X"41",  -- 65
        63333 => X"39",  -- 57
        63334 => X"36",  -- 54
        63335 => X"39",  -- 57
        63336 => X"3D",  -- 61
        63337 => X"3D",  -- 61
        63338 => X"3E",  -- 62
        63339 => X"3F",  -- 63
        63340 => X"41",  -- 65
        63341 => X"44",  -- 68
        63342 => X"45",  -- 69
        63343 => X"45",  -- 69
        63344 => X"44",  -- 68
        63345 => X"3F",  -- 63
        63346 => X"43",  -- 67
        63347 => X"49",  -- 73
        63348 => X"4C",  -- 76
        63349 => X"58",  -- 88
        63350 => X"62",  -- 98
        63351 => X"5E",  -- 94
        63352 => X"59",  -- 89
        63353 => X"4D",  -- 77
        63354 => X"47",  -- 71
        63355 => X"4E",  -- 78
        63356 => X"56",  -- 86
        63357 => X"59",  -- 89
        63358 => X"5A",  -- 90
        63359 => X"5C",  -- 92
        63360 => X"70",  -- 112
        63361 => X"71",  -- 113
        63362 => X"73",  -- 115
        63363 => X"73",  -- 115
        63364 => X"73",  -- 115
        63365 => X"73",  -- 115
        63366 => X"74",  -- 116
        63367 => X"75",  -- 117
        63368 => X"78",  -- 120
        63369 => X"70",  -- 112
        63370 => X"68",  -- 104
        63371 => X"65",  -- 101
        63372 => X"64",  -- 100
        63373 => X"66",  -- 102
        63374 => X"6F",  -- 111
        63375 => X"78",  -- 120
        63376 => X"67",  -- 103
        63377 => X"65",  -- 101
        63378 => X"66",  -- 102
        63379 => X"5F",  -- 95
        63380 => X"59",  -- 89
        63381 => X"69",  -- 105
        63382 => X"70",  -- 112
        63383 => X"5C",  -- 92
        63384 => X"74",  -- 116
        63385 => X"92",  -- 146
        63386 => X"6A",  -- 106
        63387 => X"59",  -- 89
        63388 => X"5F",  -- 95
        63389 => X"58",  -- 88
        63390 => X"76",  -- 118
        63391 => X"8D",  -- 141
        63392 => X"6F",  -- 111
        63393 => X"49",  -- 73
        63394 => X"8B",  -- 139
        63395 => X"51",  -- 81
        63396 => X"56",  -- 86
        63397 => X"59",  -- 89
        63398 => X"5A",  -- 90
        63399 => X"4E",  -- 78
        63400 => X"55",  -- 85
        63401 => X"7F",  -- 127
        63402 => X"52",  -- 82
        63403 => X"83",  -- 131
        63404 => X"8A",  -- 138
        63405 => X"39",  -- 57
        63406 => X"57",  -- 87
        63407 => X"6E",  -- 110
        63408 => X"60",  -- 96
        63409 => X"3F",  -- 63
        63410 => X"7E",  -- 126
        63411 => X"7D",  -- 125
        63412 => X"5F",  -- 95
        63413 => X"8D",  -- 141
        63414 => X"6A",  -- 106
        63415 => X"64",  -- 100
        63416 => X"67",  -- 103
        63417 => X"65",  -- 101
        63418 => X"74",  -- 116
        63419 => X"58",  -- 88
        63420 => X"84",  -- 132
        63421 => X"61",  -- 97
        63422 => X"44",  -- 68
        63423 => X"41",  -- 65
        63424 => X"57",  -- 87
        63425 => X"6C",  -- 108
        63426 => X"41",  -- 65
        63427 => X"53",  -- 83
        63428 => X"65",  -- 101
        63429 => X"46",  -- 70
        63430 => X"3A",  -- 58
        63431 => X"48",  -- 72
        63432 => X"45",  -- 69
        63433 => X"43",  -- 67
        63434 => X"4F",  -- 79
        63435 => X"57",  -- 87
        63436 => X"5B",  -- 91
        63437 => X"62",  -- 98
        63438 => X"70",  -- 112
        63439 => X"63",  -- 99
        63440 => X"5F",  -- 95
        63441 => X"67",  -- 103
        63442 => X"74",  -- 116
        63443 => X"67",  -- 103
        63444 => X"57",  -- 87
        63445 => X"50",  -- 80
        63446 => X"46",  -- 70
        63447 => X"4A",  -- 74
        63448 => X"62",  -- 98
        63449 => X"53",  -- 83
        63450 => X"43",  -- 67
        63451 => X"42",  -- 66
        63452 => X"4C",  -- 76
        63453 => X"4F",  -- 79
        63454 => X"45",  -- 69
        63455 => X"3B",  -- 59
        63456 => X"53",  -- 83
        63457 => X"61",  -- 97
        63458 => X"2E",  -- 46
        63459 => X"49",  -- 73
        63460 => X"61",  -- 97
        63461 => X"6D",  -- 109
        63462 => X"5E",  -- 94
        63463 => X"68",  -- 104
        63464 => X"5C",  -- 92
        63465 => X"5B",  -- 91
        63466 => X"7F",  -- 127
        63467 => X"78",  -- 120
        63468 => X"71",  -- 113
        63469 => X"79",  -- 121
        63470 => X"81",  -- 129
        63471 => X"7B",  -- 123
        63472 => X"7E",  -- 126
        63473 => X"71",  -- 113
        63474 => X"6D",  -- 109
        63475 => X"6A",  -- 106
        63476 => X"6F",  -- 111
        63477 => X"51",  -- 81
        63478 => X"42",  -- 66
        63479 => X"60",  -- 96
        63480 => X"4C",  -- 76
        63481 => X"5A",  -- 90
        63482 => X"45",  -- 69
        63483 => X"68",  -- 104
        63484 => X"61",  -- 97
        63485 => X"53",  -- 83
        63486 => X"53",  -- 83
        63487 => X"57",  -- 87
        63488 => X"63",  -- 99
        63489 => X"6D",  -- 109
        63490 => X"5E",  -- 94
        63491 => X"4E",  -- 78
        63492 => X"48",  -- 72
        63493 => X"74",  -- 116
        63494 => X"7E",  -- 126
        63495 => X"78",  -- 120
        63496 => X"43",  -- 67
        63497 => X"3F",  -- 63
        63498 => X"53",  -- 83
        63499 => X"96",  -- 150
        63500 => X"69",  -- 105
        63501 => X"54",  -- 84
        63502 => X"33",  -- 51
        63503 => X"72",  -- 114
        63504 => X"5E",  -- 94
        63505 => X"76",  -- 118
        63506 => X"83",  -- 131
        63507 => X"43",  -- 67
        63508 => X"51",  -- 81
        63509 => X"57",  -- 87
        63510 => X"4A",  -- 74
        63511 => X"4B",  -- 75
        63512 => X"49",  -- 73
        63513 => X"92",  -- 146
        63514 => X"51",  -- 81
        63515 => X"78",  -- 120
        63516 => X"51",  -- 81
        63517 => X"7B",  -- 123
        63518 => X"45",  -- 69
        63519 => X"2A",  -- 42
        63520 => X"15",  -- 21
        63521 => X"11",  -- 17
        63522 => X"10",  -- 16
        63523 => X"16",  -- 22
        63524 => X"19",  -- 25
        63525 => X"17",  -- 23
        63526 => X"19",  -- 25
        63527 => X"1A",  -- 26
        63528 => X"20",  -- 32
        63529 => X"1F",  -- 31
        63530 => X"1C",  -- 28
        63531 => X"28",  -- 40
        63532 => X"1E",  -- 30
        63533 => X"21",  -- 33
        63534 => X"28",  -- 40
        63535 => X"65",  -- 101
        63536 => X"25",  -- 37
        63537 => X"20",  -- 32
        63538 => X"1D",  -- 29
        63539 => X"1C",  -- 28
        63540 => X"1D",  -- 29
        63541 => X"1F",  -- 31
        63542 => X"20",  -- 32
        63543 => X"20",  -- 32
        63544 => X"23",  -- 35
        63545 => X"25",  -- 37
        63546 => X"24",  -- 36
        63547 => X"27",  -- 39
        63548 => X"2F",  -- 47
        63549 => X"38",  -- 56
        63550 => X"3A",  -- 58
        63551 => X"36",  -- 54
        63552 => X"2C",  -- 44
        63553 => X"30",  -- 48
        63554 => X"3F",  -- 63
        63555 => X"51",  -- 81
        63556 => X"5B",  -- 91
        63557 => X"5A",  -- 90
        63558 => X"5F",  -- 95
        63559 => X"68",  -- 104
        63560 => X"6A",  -- 106
        63561 => X"5F",  -- 95
        63562 => X"4C",  -- 76
        63563 => X"39",  -- 57
        63564 => X"2F",  -- 47
        63565 => X"2F",  -- 47
        63566 => X"31",  -- 49
        63567 => X"30",  -- 48
        63568 => X"43",  -- 67
        63569 => X"64",  -- 100
        63570 => X"45",  -- 69
        63571 => X"6A",  -- 106
        63572 => X"8E",  -- 142
        63573 => X"7C",  -- 124
        63574 => X"77",  -- 119
        63575 => X"71",  -- 113
        63576 => X"76",  -- 118
        63577 => X"6F",  -- 111
        63578 => X"69",  -- 105
        63579 => X"67",  -- 103
        63580 => X"70",  -- 112
        63581 => X"5B",  -- 91
        63582 => X"2E",  -- 46
        63583 => X"26",  -- 38
        63584 => X"3E",  -- 62
        63585 => X"8C",  -- 140
        63586 => X"B1",  -- 177
        63587 => X"93",  -- 147
        63588 => X"B5",  -- 181
        63589 => X"A7",  -- 167
        63590 => X"AE",  -- 174
        63591 => X"8F",  -- 143
        63592 => X"A6",  -- 166
        63593 => X"93",  -- 147
        63594 => X"9C",  -- 156
        63595 => X"4F",  -- 79
        63596 => X"04",  -- 4
        63597 => X"06",  -- 6
        63598 => X"09",  -- 9
        63599 => X"0C",  -- 12
        63600 => X"59",  -- 89
        63601 => X"89",  -- 137
        63602 => X"95",  -- 149
        63603 => X"6E",  -- 110
        63604 => X"2C",  -- 44
        63605 => X"39",  -- 57
        63606 => X"8C",  -- 140
        63607 => X"C1",  -- 193
        63608 => X"C1",  -- 193
        63609 => X"C1",  -- 193
        63610 => X"B7",  -- 183
        63611 => X"B1",  -- 177
        63612 => X"BB",  -- 187
        63613 => X"C1",  -- 193
        63614 => X"C0",  -- 192
        63615 => X"C2",  -- 194
        63616 => X"C4",  -- 196
        63617 => X"BB",  -- 187
        63618 => X"B3",  -- 179
        63619 => X"B8",  -- 184
        63620 => X"C9",  -- 201
        63621 => X"B0",  -- 176
        63622 => X"84",  -- 132
        63623 => X"80",  -- 128
        63624 => X"B5",  -- 181
        63625 => X"C2",  -- 194
        63626 => X"C5",  -- 197
        63627 => X"B9",  -- 185
        63628 => X"B6",  -- 182
        63629 => X"C0",  -- 192
        63630 => X"C9",  -- 201
        63631 => X"C7",  -- 199
        63632 => X"CB",  -- 203
        63633 => X"CF",  -- 207
        63634 => X"CA",  -- 202
        63635 => X"CA",  -- 202
        63636 => X"9C",  -- 156
        63637 => X"52",  -- 82
        63638 => X"3D",  -- 61
        63639 => X"40",  -- 64
        63640 => X"38",  -- 56
        63641 => X"2F",  -- 47
        63642 => X"2B",  -- 43
        63643 => X"31",  -- 49
        63644 => X"3D",  -- 61
        63645 => X"44",  -- 68
        63646 => X"49",  -- 73
        63647 => X"4C",  -- 76
        63648 => X"50",  -- 80
        63649 => X"5B",  -- 91
        63650 => X"61",  -- 97
        63651 => X"5C",  -- 92
        63652 => X"4D",  -- 77
        63653 => X"41",  -- 65
        63654 => X"3D",  -- 61
        63655 => X"3F",  -- 63
        63656 => X"42",  -- 66
        63657 => X"3D",  -- 61
        63658 => X"37",  -- 55
        63659 => X"37",  -- 55
        63660 => X"39",  -- 57
        63661 => X"3C",  -- 60
        63662 => X"3D",  -- 61
        63663 => X"3D",  -- 61
        63664 => X"3D",  -- 61
        63665 => X"38",  -- 56
        63666 => X"3E",  -- 62
        63667 => X"45",  -- 69
        63668 => X"47",  -- 71
        63669 => X"4D",  -- 77
        63670 => X"51",  -- 81
        63671 => X"4E",  -- 78
        63672 => X"4E",  -- 78
        63673 => X"44",  -- 68
        63674 => X"41",  -- 65
        63675 => X"44",  -- 68
        63676 => X"49",  -- 73
        63677 => X"52",  -- 82
        63678 => X"58",  -- 88
        63679 => X"55",  -- 85
        63680 => X"6C",  -- 108
        63681 => X"6D",  -- 109
        63682 => X"6E",  -- 110
        63683 => X"6F",  -- 111
        63684 => X"70",  -- 112
        63685 => X"73",  -- 115
        63686 => X"77",  -- 119
        63687 => X"7A",  -- 122
        63688 => X"72",  -- 114
        63689 => X"6C",  -- 108
        63690 => X"69",  -- 105
        63691 => X"6C",  -- 108
        63692 => X"6E",  -- 110
        63693 => X"6D",  -- 109
        63694 => X"6D",  -- 109
        63695 => X"70",  -- 112
        63696 => X"77",  -- 119
        63697 => X"6F",  -- 111
        63698 => X"68",  -- 104
        63699 => X"6B",  -- 107
        63700 => X"6B",  -- 107
        63701 => X"61",  -- 97
        63702 => X"60",  -- 96
        63703 => X"6E",  -- 110
        63704 => X"82",  -- 130
        63705 => X"6A",  -- 106
        63706 => X"5A",  -- 90
        63707 => X"58",  -- 88
        63708 => X"61",  -- 97
        63709 => X"75",  -- 117
        63710 => X"75",  -- 117
        63711 => X"5B",  -- 91
        63712 => X"4A",  -- 74
        63713 => X"63",  -- 99
        63714 => X"66",  -- 102
        63715 => X"50",  -- 80
        63716 => X"58",  -- 88
        63717 => X"63",  -- 99
        63718 => X"53",  -- 83
        63719 => X"58",  -- 88
        63720 => X"68",  -- 104
        63721 => X"70",  -- 112
        63722 => X"6F",  -- 111
        63723 => X"AD",  -- 173
        63724 => X"4C",  -- 76
        63725 => X"59",  -- 89
        63726 => X"63",  -- 99
        63727 => X"6F",  -- 111
        63728 => X"42",  -- 66
        63729 => X"60",  -- 96
        63730 => X"78",  -- 120
        63731 => X"67",  -- 103
        63732 => X"70",  -- 112
        63733 => X"83",  -- 131
        63734 => X"4B",  -- 75
        63735 => X"79",  -- 121
        63736 => X"5E",  -- 94
        63737 => X"6C",  -- 108
        63738 => X"69",  -- 105
        63739 => X"66",  -- 102
        63740 => X"7C",  -- 124
        63741 => X"54",  -- 84
        63742 => X"40",  -- 64
        63743 => X"56",  -- 86
        63744 => X"70",  -- 112
        63745 => X"3F",  -- 63
        63746 => X"58",  -- 88
        63747 => X"5A",  -- 90
        63748 => X"65",  -- 101
        63749 => X"39",  -- 57
        63750 => X"51",  -- 81
        63751 => X"48",  -- 72
        63752 => X"42",  -- 66
        63753 => X"44",  -- 68
        63754 => X"4F",  -- 79
        63755 => X"5C",  -- 92
        63756 => X"58",  -- 88
        63757 => X"68",  -- 104
        63758 => X"72",  -- 114
        63759 => X"59",  -- 89
        63760 => X"6E",  -- 110
        63761 => X"75",  -- 117
        63762 => X"74",  -- 116
        63763 => X"5D",  -- 93
        63764 => X"65",  -- 101
        63765 => X"7F",  -- 127
        63766 => X"70",  -- 112
        63767 => X"56",  -- 86
        63768 => X"6E",  -- 110
        63769 => X"47",  -- 71
        63770 => X"3E",  -- 62
        63771 => X"57",  -- 87
        63772 => X"64",  -- 100
        63773 => X"5B",  -- 91
        63774 => X"53",  -- 83
        63775 => X"53",  -- 83
        63776 => X"5A",  -- 90
        63777 => X"7F",  -- 127
        63778 => X"46",  -- 70
        63779 => X"50",  -- 80
        63780 => X"65",  -- 101
        63781 => X"74",  -- 116
        63782 => X"61",  -- 97
        63783 => X"6D",  -- 109
        63784 => X"7B",  -- 123
        63785 => X"5B",  -- 91
        63786 => X"77",  -- 119
        63787 => X"99",  -- 153
        63788 => X"7D",  -- 125
        63789 => X"7E",  -- 126
        63790 => X"79",  -- 121
        63791 => X"87",  -- 135
        63792 => X"84",  -- 132
        63793 => X"79",  -- 121
        63794 => X"72",  -- 114
        63795 => X"73",  -- 115
        63796 => X"6B",  -- 107
        63797 => X"77",  -- 119
        63798 => X"50",  -- 80
        63799 => X"50",  -- 80
        63800 => X"51",  -- 81
        63801 => X"55",  -- 85
        63802 => X"52",  -- 82
        63803 => X"59",  -- 89
        63804 => X"6D",  -- 109
        63805 => X"51",  -- 81
        63806 => X"59",  -- 89
        63807 => X"4B",  -- 75
        63808 => X"52",  -- 82
        63809 => X"6C",  -- 108
        63810 => X"56",  -- 86
        63811 => X"5A",  -- 90
        63812 => X"4F",  -- 79
        63813 => X"67",  -- 103
        63814 => X"71",  -- 113
        63815 => X"7E",  -- 126
        63816 => X"6B",  -- 107
        63817 => X"50",  -- 80
        63818 => X"4D",  -- 77
        63819 => X"66",  -- 102
        63820 => X"92",  -- 146
        63821 => X"5E",  -- 94
        63822 => X"55",  -- 85
        63823 => X"47",  -- 71
        63824 => X"80",  -- 128
        63825 => X"5B",  -- 91
        63826 => X"B0",  -- 176
        63827 => X"64",  -- 100
        63828 => X"43",  -- 67
        63829 => X"61",  -- 97
        63830 => X"4B",  -- 75
        63831 => X"48",  -- 72
        63832 => X"4B",  -- 75
        63833 => X"52",  -- 82
        63834 => X"87",  -- 135
        63835 => X"5B",  -- 91
        63836 => X"5A",  -- 90
        63837 => X"45",  -- 69
        63838 => X"6D",  -- 109
        63839 => X"13",  -- 19
        63840 => X"0E",  -- 14
        63841 => X"10",  -- 16
        63842 => X"13",  -- 19
        63843 => X"16",  -- 22
        63844 => X"18",  -- 24
        63845 => X"1A",  -- 26
        63846 => X"1C",  -- 28
        63847 => X"1E",  -- 30
        63848 => X"20",  -- 32
        63849 => X"29",  -- 41
        63850 => X"2D",  -- 45
        63851 => X"1A",  -- 26
        63852 => X"21",  -- 33
        63853 => X"18",  -- 24
        63854 => X"0B",  -- 11
        63855 => X"24",  -- 36
        63856 => X"26",  -- 38
        63857 => X"1F",  -- 31
        63858 => X"17",  -- 23
        63859 => X"16",  -- 22
        63860 => X"1B",  -- 27
        63861 => X"1E",  -- 30
        63862 => X"22",  -- 34
        63863 => X"22",  -- 34
        63864 => X"2D",  -- 45
        63865 => X"32",  -- 50
        63866 => X"32",  -- 50
        63867 => X"32",  -- 50
        63868 => X"35",  -- 53
        63869 => X"3A",  -- 58
        63870 => X"3C",  -- 60
        63871 => X"39",  -- 57
        63872 => X"2E",  -- 46
        63873 => X"31",  -- 49
        63874 => X"3B",  -- 59
        63875 => X"4E",  -- 78
        63876 => X"5B",  -- 91
        63877 => X"63",  -- 99
        63878 => X"6F",  -- 111
        63879 => X"7D",  -- 125
        63880 => X"75",  -- 117
        63881 => X"67",  -- 103
        63882 => X"4E",  -- 78
        63883 => X"39",  -- 57
        63884 => X"2F",  -- 47
        63885 => X"2F",  -- 47
        63886 => X"2E",  -- 46
        63887 => X"2B",  -- 43
        63888 => X"3B",  -- 59
        63889 => X"53",  -- 83
        63890 => X"4B",  -- 75
        63891 => X"77",  -- 119
        63892 => X"76",  -- 118
        63893 => X"6A",  -- 106
        63894 => X"6C",  -- 108
        63895 => X"68",  -- 104
        63896 => X"74",  -- 116
        63897 => X"69",  -- 105
        63898 => X"6D",  -- 109
        63899 => X"6D",  -- 109
        63900 => X"6F",  -- 111
        63901 => X"65",  -- 101
        63902 => X"45",  -- 69
        63903 => X"37",  -- 55
        63904 => X"63",  -- 99
        63905 => X"97",  -- 151
        63906 => X"92",  -- 146
        63907 => X"A8",  -- 168
        63908 => X"AF",  -- 175
        63909 => X"A5",  -- 165
        63910 => X"92",  -- 146
        63911 => X"97",  -- 151
        63912 => X"A4",  -- 164
        63913 => X"A7",  -- 167
        63914 => X"8F",  -- 143
        63915 => X"5E",  -- 94
        63916 => X"00",  -- 0
        63917 => X"05",  -- 5
        63918 => X"02",  -- 2
        63919 => X"05",  -- 5
        63920 => X"32",  -- 50
        63921 => X"81",  -- 129
        63922 => X"98",  -- 152
        63923 => X"89",  -- 137
        63924 => X"59",  -- 89
        63925 => X"36",  -- 54
        63926 => X"7A",  -- 122
        63927 => X"C2",  -- 194
        63928 => X"C5",  -- 197
        63929 => X"C0",  -- 192
        63930 => X"B0",  -- 176
        63931 => X"A7",  -- 167
        63932 => X"AE",  -- 174
        63933 => X"B5",  -- 181
        63934 => X"B5",  -- 181
        63935 => X"B8",  -- 184
        63936 => X"BB",  -- 187
        63937 => X"B6",  -- 182
        63938 => X"B4",  -- 180
        63939 => X"AC",  -- 172
        63940 => X"C3",  -- 195
        63941 => X"BF",  -- 191
        63942 => X"7C",  -- 124
        63943 => X"5B",  -- 91
        63944 => X"AA",  -- 170
        63945 => X"C3",  -- 195
        63946 => X"C2",  -- 194
        63947 => X"A2",  -- 162
        63948 => X"97",  -- 151
        63949 => X"B1",  -- 177
        63950 => X"C6",  -- 198
        63951 => X"C5",  -- 197
        63952 => X"CE",  -- 206
        63953 => X"D3",  -- 211
        63954 => X"CD",  -- 205
        63955 => X"C8",  -- 200
        63956 => X"91",  -- 145
        63957 => X"47",  -- 71
        63958 => X"3C",  -- 60
        63959 => X"41",  -- 65
        63960 => X"34",  -- 52
        63961 => X"2B",  -- 43
        63962 => X"26",  -- 38
        63963 => X"2D",  -- 45
        63964 => X"38",  -- 56
        63965 => X"43",  -- 67
        63966 => X"4B",  -- 75
        63967 => X"4E",  -- 78
        63968 => X"5B",  -- 91
        63969 => X"64",  -- 100
        63970 => X"6A",  -- 106
        63971 => X"64",  -- 100
        63972 => X"54",  -- 84
        63973 => X"44",  -- 68
        63974 => X"40",  -- 64
        63975 => X"42",  -- 66
        63976 => X"47",  -- 71
        63977 => X"3B",  -- 59
        63978 => X"31",  -- 49
        63979 => X"2C",  -- 44
        63980 => X"32",  -- 50
        63981 => X"37",  -- 55
        63982 => X"38",  -- 56
        63983 => X"35",  -- 53
        63984 => X"3C",  -- 60
        63985 => X"37",  -- 55
        63986 => X"3C",  -- 60
        63987 => X"44",  -- 68
        63988 => X"43",  -- 67
        63989 => X"45",  -- 69
        63990 => X"49",  -- 73
        63991 => X"45",  -- 69
        63992 => X"47",  -- 71
        63993 => X"40",  -- 64
        63994 => X"3D",  -- 61
        63995 => X"3C",  -- 60
        63996 => X"41",  -- 65
        63997 => X"4E",  -- 78
        63998 => X"56",  -- 86
        63999 => X"50",  -- 80
        64000 => X"6E",  -- 110
        64001 => X"70",  -- 112
        64002 => X"68",  -- 104
        64003 => X"6C",  -- 108
        64004 => X"79",  -- 121
        64005 => X"74",  -- 116
        64006 => X"70",  -- 112
        64007 => X"80",  -- 128
        64008 => X"6C",  -- 108
        64009 => X"72",  -- 114
        64010 => X"73",  -- 115
        64011 => X"6D",  -- 109
        64012 => X"6C",  -- 108
        64013 => X"72",  -- 114
        64014 => X"74",  -- 116
        64015 => X"71",  -- 113
        64016 => X"6F",  -- 111
        64017 => X"64",  -- 100
        64018 => X"73",  -- 115
        64019 => X"6A",  -- 106
        64020 => X"61",  -- 97
        64021 => X"66",  -- 102
        64022 => X"63",  -- 99
        64023 => X"79",  -- 121
        64024 => X"7B",  -- 123
        64025 => X"4F",  -- 79
        64026 => X"45",  -- 69
        64027 => X"55",  -- 85
        64028 => X"6B",  -- 107
        64029 => X"84",  -- 132
        64030 => X"5C",  -- 92
        64031 => X"6A",  -- 106
        64032 => X"46",  -- 70
        64033 => X"67",  -- 103
        64034 => X"4C",  -- 76
        64035 => X"4E",  -- 78
        64036 => X"4F",  -- 79
        64037 => X"5B",  -- 91
        64038 => X"5A",  -- 90
        64039 => X"5A",  -- 90
        64040 => X"7C",  -- 124
        64041 => X"5F",  -- 95
        64042 => X"9D",  -- 157
        64043 => X"75",  -- 117
        64044 => X"4C",  -- 76
        64045 => X"5B",  -- 91
        64046 => X"85",  -- 133
        64047 => X"52",  -- 82
        64048 => X"56",  -- 86
        64049 => X"74",  -- 116
        64050 => X"78",  -- 120
        64051 => X"54",  -- 84
        64052 => X"91",  -- 145
        64053 => X"51",  -- 81
        64054 => X"6E",  -- 110
        64055 => X"69",  -- 105
        64056 => X"6D",  -- 109
        64057 => X"6E",  -- 110
        64058 => X"57",  -- 87
        64059 => X"85",  -- 133
        64060 => X"49",  -- 73
        64061 => X"32",  -- 50
        64062 => X"53",  -- 83
        64063 => X"65",  -- 101
        64064 => X"3D",  -- 61
        64065 => X"3D",  -- 61
        64066 => X"49",  -- 73
        64067 => X"57",  -- 87
        64068 => X"4E",  -- 78
        64069 => X"36",  -- 54
        64070 => X"2E",  -- 46
        64071 => X"36",  -- 54
        64072 => X"2C",  -- 44
        64073 => X"31",  -- 49
        64074 => X"46",  -- 70
        64075 => X"76",  -- 118
        64076 => X"65",  -- 101
        64077 => X"64",  -- 100
        64078 => X"6E",  -- 110
        64079 => X"6D",  -- 109
        64080 => X"65",  -- 101
        64081 => X"81",  -- 129
        64082 => X"71",  -- 113
        64083 => X"84",  -- 132
        64084 => X"70",  -- 112
        64085 => X"69",  -- 105
        64086 => X"7A",  -- 122
        64087 => X"79",  -- 121
        64088 => X"6F",  -- 111
        64089 => X"51",  -- 81
        64090 => X"4B",  -- 75
        64091 => X"82",  -- 130
        64092 => X"62",  -- 98
        64093 => X"4D",  -- 77
        64094 => X"5E",  -- 94
        64095 => X"67",  -- 103
        64096 => X"6F",  -- 111
        64097 => X"51",  -- 81
        64098 => X"6B",  -- 107
        64099 => X"83",  -- 131
        64100 => X"54",  -- 84
        64101 => X"6F",  -- 111
        64102 => X"65",  -- 101
        64103 => X"7E",  -- 126
        64104 => X"70",  -- 112
        64105 => X"7C",  -- 124
        64106 => X"86",  -- 134
        64107 => X"9D",  -- 157
        64108 => X"96",  -- 150
        64109 => X"86",  -- 134
        64110 => X"99",  -- 153
        64111 => X"9A",  -- 154
        64112 => X"79",  -- 121
        64113 => X"88",  -- 136
        64114 => X"88",  -- 136
        64115 => X"72",  -- 114
        64116 => X"76",  -- 118
        64117 => X"76",  -- 118
        64118 => X"4D",  -- 77
        64119 => X"49",  -- 73
        64120 => X"47",  -- 71
        64121 => X"57",  -- 87
        64122 => X"45",  -- 69
        64123 => X"4A",  -- 74
        64124 => X"5F",  -- 95
        64125 => X"6D",  -- 109
        64126 => X"45",  -- 69
        64127 => X"4A",  -- 74
        64128 => X"4D",  -- 77
        64129 => X"6B",  -- 107
        64130 => X"71",  -- 113
        64131 => X"58",  -- 88
        64132 => X"5B",  -- 91
        64133 => X"6B",  -- 107
        64134 => X"65",  -- 101
        64135 => X"6C",  -- 108
        64136 => X"89",  -- 137
        64137 => X"6C",  -- 108
        64138 => X"4E",  -- 78
        64139 => X"63",  -- 99
        64140 => X"63",  -- 99
        64141 => X"9A",  -- 154
        64142 => X"5C",  -- 92
        64143 => X"41",  -- 65
        64144 => X"73",  -- 115
        64145 => X"5F",  -- 95
        64146 => X"87",  -- 135
        64147 => X"97",  -- 151
        64148 => X"4B",  -- 75
        64149 => X"4D",  -- 77
        64150 => X"56",  -- 86
        64151 => X"47",  -- 71
        64152 => X"42",  -- 66
        64153 => X"41",  -- 65
        64154 => X"5E",  -- 94
        64155 => X"56",  -- 86
        64156 => X"48",  -- 72
        64157 => X"55",  -- 85
        64158 => X"30",  -- 48
        64159 => X"57",  -- 87
        64160 => X"01",  -- 1
        64161 => X"16",  -- 22
        64162 => X"17",  -- 23
        64163 => X"09",  -- 9
        64164 => X"19",  -- 25
        64165 => X"29",  -- 41
        64166 => X"1D",  -- 29
        64167 => X"1D",  -- 29
        64168 => X"19",  -- 25
        64169 => X"1D",  -- 29
        64170 => X"26",  -- 38
        64171 => X"2C",  -- 44
        64172 => X"29",  -- 41
        64173 => X"20",  -- 32
        64174 => X"1A",  -- 26
        64175 => X"19",  -- 25
        64176 => X"16",  -- 22
        64177 => X"16",  -- 22
        64178 => X"17",  -- 23
        64179 => X"1B",  -- 27
        64180 => X"1C",  -- 28
        64181 => X"20",  -- 32
        64182 => X"23",  -- 35
        64183 => X"26",  -- 38
        64184 => X"25",  -- 37
        64185 => X"2B",  -- 43
        64186 => X"2F",  -- 47
        64187 => X"33",  -- 51
        64188 => X"37",  -- 55
        64189 => X"3E",  -- 62
        64190 => X"40",  -- 64
        64191 => X"3F",  -- 63
        64192 => X"32",  -- 50
        64193 => X"32",  -- 50
        64194 => X"36",  -- 54
        64195 => X"44",  -- 68
        64196 => X"59",  -- 89
        64197 => X"6E",  -- 110
        64198 => X"82",  -- 130
        64199 => X"91",  -- 145
        64200 => X"8C",  -- 140
        64201 => X"70",  -- 112
        64202 => X"49",  -- 73
        64203 => X"2E",  -- 46
        64204 => X"2A",  -- 42
        64205 => X"31",  -- 49
        64206 => X"33",  -- 51
        64207 => X"2F",  -- 47
        64208 => X"43",  -- 67
        64209 => X"43",  -- 67
        64210 => X"5B",  -- 91
        64211 => X"72",  -- 114
        64212 => X"82",  -- 130
        64213 => X"7A",  -- 122
        64214 => X"68",  -- 104
        64215 => X"71",  -- 113
        64216 => X"6E",  -- 110
        64217 => X"6B",  -- 107
        64218 => X"6F",  -- 111
        64219 => X"6D",  -- 109
        64220 => X"74",  -- 116
        64221 => X"71",  -- 113
        64222 => X"5F",  -- 95
        64223 => X"61",  -- 97
        64224 => X"87",  -- 135
        64225 => X"83",  -- 131
        64226 => X"92",  -- 146
        64227 => X"9E",  -- 158
        64228 => X"93",  -- 147
        64229 => X"89",  -- 137
        64230 => X"8E",  -- 142
        64231 => X"98",  -- 152
        64232 => X"9F",  -- 159
        64233 => X"B1",  -- 177
        64234 => X"6A",  -- 106
        64235 => X"40",  -- 64
        64236 => X"10",  -- 16
        64237 => X"00",  -- 0
        64238 => X"03",  -- 3
        64239 => X"08",  -- 8
        64240 => X"23",  -- 35
        64241 => X"57",  -- 87
        64242 => X"92",  -- 146
        64243 => X"93",  -- 147
        64244 => X"93",  -- 147
        64245 => X"6D",  -- 109
        64246 => X"98",  -- 152
        64247 => X"BA",  -- 186
        64248 => X"CE",  -- 206
        64249 => X"B1",  -- 177
        64250 => X"A3",  -- 163
        64251 => X"9B",  -- 155
        64252 => X"A9",  -- 169
        64253 => X"A4",  -- 164
        64254 => X"B4",  -- 180
        64255 => X"BA",  -- 186
        64256 => X"B9",  -- 185
        64257 => X"AD",  -- 173
        64258 => X"B9",  -- 185
        64259 => X"B0",  -- 176
        64260 => X"AA",  -- 170
        64261 => X"BC",  -- 188
        64262 => X"9C",  -- 156
        64263 => X"5D",  -- 93
        64264 => X"94",  -- 148
        64265 => X"CE",  -- 206
        64266 => X"BC",  -- 188
        64267 => X"7F",  -- 127
        64268 => X"97",  -- 151
        64269 => X"A2",  -- 162
        64270 => X"B3",  -- 179
        64271 => X"D6",  -- 214
        64272 => X"D9",  -- 217
        64273 => X"D0",  -- 208
        64274 => X"D3",  -- 211
        64275 => X"BA",  -- 186
        64276 => X"79",  -- 121
        64277 => X"45",  -- 69
        64278 => X"3A",  -- 58
        64279 => X"3B",  -- 59
        64280 => X"35",  -- 53
        64281 => X"30",  -- 48
        64282 => X"22",  -- 34
        64283 => X"28",  -- 40
        64284 => X"3D",  -- 61
        64285 => X"42",  -- 66
        64286 => X"42",  -- 66
        64287 => X"53",  -- 83
        64288 => X"5C",  -- 92
        64289 => X"67",  -- 103
        64290 => X"6E",  -- 110
        64291 => X"67",  -- 103
        64292 => X"53",  -- 83
        64293 => X"44",  -- 68
        64294 => X"42",  -- 66
        64295 => X"48",  -- 72
        64296 => X"47",  -- 71
        64297 => X"43",  -- 67
        64298 => X"38",  -- 56
        64299 => X"2B",  -- 43
        64300 => X"27",  -- 39
        64301 => X"2C",  -- 44
        64302 => X"31",  -- 49
        64303 => X"32",  -- 50
        64304 => X"39",  -- 57
        64305 => X"31",  -- 49
        64306 => X"3E",  -- 62
        64307 => X"3A",  -- 58
        64308 => X"43",  -- 67
        64309 => X"3C",  -- 60
        64310 => X"46",  -- 70
        64311 => X"3C",  -- 60
        64312 => X"3E",  -- 62
        64313 => X"3D",  -- 61
        64314 => X"3A",  -- 58
        64315 => X"36",  -- 54
        64316 => X"3C",  -- 60
        64317 => X"47",  -- 71
        64318 => X"4B",  -- 75
        64319 => X"4A",  -- 74
        64320 => X"75",  -- 117
        64321 => X"74",  -- 116
        64322 => X"6B",  -- 107
        64323 => X"6D",  -- 109
        64324 => X"76",  -- 118
        64325 => X"6C",  -- 108
        64326 => X"63",  -- 99
        64327 => X"6C",  -- 108
        64328 => X"71",  -- 113
        64329 => X"71",  -- 113
        64330 => X"6D",  -- 109
        64331 => X"69",  -- 105
        64332 => X"68",  -- 104
        64333 => X"6C",  -- 108
        64334 => X"6E",  -- 110
        64335 => X"6E",  -- 110
        64336 => X"69",  -- 105
        64337 => X"72",  -- 114
        64338 => X"67",  -- 103
        64339 => X"6F",  -- 111
        64340 => X"6A",  -- 106
        64341 => X"62",  -- 98
        64342 => X"66",  -- 102
        64343 => X"87",  -- 135
        64344 => X"58",  -- 88
        64345 => X"55",  -- 85
        64346 => X"5C",  -- 92
        64347 => X"5B",  -- 91
        64348 => X"69",  -- 105
        64349 => X"70",  -- 112
        64350 => X"64",  -- 100
        64351 => X"56",  -- 86
        64352 => X"4C",  -- 76
        64353 => X"58",  -- 88
        64354 => X"38",  -- 56
        64355 => X"33",  -- 51
        64356 => X"3B",  -- 59
        64357 => X"44",  -- 68
        64358 => X"43",  -- 67
        64359 => X"77",  -- 119
        64360 => X"7E",  -- 126
        64361 => X"87",  -- 135
        64362 => X"85",  -- 133
        64363 => X"51",  -- 81
        64364 => X"51",  -- 81
        64365 => X"7C",  -- 124
        64366 => X"63",  -- 99
        64367 => X"4D",  -- 77
        64368 => X"63",  -- 99
        64369 => X"82",  -- 130
        64370 => X"63",  -- 99
        64371 => X"7F",  -- 127
        64372 => X"53",  -- 83
        64373 => X"55",  -- 85
        64374 => X"78",  -- 120
        64375 => X"64",  -- 100
        64376 => X"58",  -- 88
        64377 => X"64",  -- 100
        64378 => X"52",  -- 82
        64379 => X"60",  -- 96
        64380 => X"3C",  -- 60
        64381 => X"47",  -- 71
        64382 => X"57",  -- 87
        64383 => X"44",  -- 68
        64384 => X"2E",  -- 46
        64385 => X"3C",  -- 60
        64386 => X"43",  -- 67
        64387 => X"3A",  -- 58
        64388 => X"2B",  -- 43
        64389 => X"21",  -- 33
        64390 => X"1C",  -- 28
        64391 => X"19",  -- 25
        64392 => X"23",  -- 35
        64393 => X"33",  -- 51
        64394 => X"4C",  -- 76
        64395 => X"6E",  -- 110
        64396 => X"65",  -- 101
        64397 => X"71",  -- 113
        64398 => X"71",  -- 113
        64399 => X"6B",  -- 107
        64400 => X"74",  -- 116
        64401 => X"86",  -- 134
        64402 => X"89",  -- 137
        64403 => X"71",  -- 113
        64404 => X"46",  -- 70
        64405 => X"68",  -- 104
        64406 => X"98",  -- 152
        64407 => X"83",  -- 131
        64408 => X"59",  -- 89
        64409 => X"5E",  -- 94
        64410 => X"6D",  -- 109
        64411 => X"7E",  -- 126
        64412 => X"5F",  -- 95
        64413 => X"52",  -- 82
        64414 => X"5D",  -- 93
        64415 => X"5F",  -- 95
        64416 => X"64",  -- 100
        64417 => X"63",  -- 99
        64418 => X"5F",  -- 95
        64419 => X"98",  -- 152
        64420 => X"81",  -- 129
        64421 => X"62",  -- 98
        64422 => X"66",  -- 102
        64423 => X"76",  -- 118
        64424 => X"92",  -- 146
        64425 => X"94",  -- 148
        64426 => X"99",  -- 153
        64427 => X"AC",  -- 172
        64428 => X"9B",  -- 155
        64429 => X"7D",  -- 125
        64430 => X"8F",  -- 143
        64431 => X"A1",  -- 161
        64432 => X"9C",  -- 156
        64433 => X"78",  -- 120
        64434 => X"7F",  -- 127
        64435 => X"7C",  -- 124
        64436 => X"5F",  -- 95
        64437 => X"66",  -- 102
        64438 => X"62",  -- 98
        64439 => X"3B",  -- 59
        64440 => X"47",  -- 71
        64441 => X"5B",  -- 91
        64442 => X"43",  -- 67
        64443 => X"4A",  -- 74
        64444 => X"52",  -- 82
        64445 => X"66",  -- 102
        64446 => X"4A",  -- 74
        64447 => X"42",  -- 66
        64448 => X"3E",  -- 62
        64449 => X"5D",  -- 93
        64450 => X"71",  -- 113
        64451 => X"52",  -- 82
        64452 => X"54",  -- 84
        64453 => X"74",  -- 116
        64454 => X"5C",  -- 92
        64455 => X"66",  -- 102
        64456 => X"73",  -- 115
        64457 => X"7D",  -- 125
        64458 => X"5A",  -- 90
        64459 => X"65",  -- 101
        64460 => X"5B",  -- 91
        64461 => X"78",  -- 120
        64462 => X"8A",  -- 138
        64463 => X"4F",  -- 79
        64464 => X"52",  -- 82
        64465 => X"7E",  -- 126
        64466 => X"55",  -- 85
        64467 => X"98",  -- 152
        64468 => X"7A",  -- 122
        64469 => X"42",  -- 66
        64470 => X"4D",  -- 77
        64471 => X"3B",  -- 59
        64472 => X"4D",  -- 77
        64473 => X"3C",  -- 60
        64474 => X"11",  -- 17
        64475 => X"6B",  -- 107
        64476 => X"2E",  -- 46
        64477 => X"43",  -- 67
        64478 => X"58",  -- 88
        64479 => X"50",  -- 80
        64480 => X"39",  -- 57
        64481 => X"04",  -- 4
        64482 => X"23",  -- 35
        64483 => X"1C",  -- 28
        64484 => X"22",  -- 34
        64485 => X"27",  -- 39
        64486 => X"1D",  -- 29
        64487 => X"32",  -- 50
        64488 => X"2B",  -- 43
        64489 => X"24",  -- 36
        64490 => X"22",  -- 34
        64491 => X"28",  -- 40
        64492 => X"2D",  -- 45
        64493 => X"2B",  -- 43
        64494 => X"25",  -- 37
        64495 => X"21",  -- 33
        64496 => X"22",  -- 34
        64497 => X"24",  -- 36
        64498 => X"27",  -- 39
        64499 => X"2A",  -- 42
        64500 => X"2D",  -- 45
        64501 => X"2C",  -- 44
        64502 => X"28",  -- 40
        64503 => X"25",  -- 37
        64504 => X"26",  -- 38
        64505 => X"2C",  -- 44
        64506 => X"31",  -- 49
        64507 => X"36",  -- 54
        64508 => X"3C",  -- 60
        64509 => X"41",  -- 65
        64510 => X"43",  -- 67
        64511 => X"41",  -- 65
        64512 => X"35",  -- 53
        64513 => X"31",  -- 49
        64514 => X"31",  -- 49
        64515 => X"40",  -- 64
        64516 => X"59",  -- 89
        64517 => X"70",  -- 112
        64518 => X"85",  -- 133
        64519 => X"91",  -- 145
        64520 => X"89",  -- 137
        64521 => X"72",  -- 114
        64522 => X"51",  -- 81
        64523 => X"3B",  -- 59
        64524 => X"38",  -- 56
        64525 => X"40",  -- 64
        64526 => X"3F",  -- 63
        64527 => X"3A",  -- 58
        64528 => X"44",  -- 68
        64529 => X"4E",  -- 78
        64530 => X"63",  -- 99
        64531 => X"6E",  -- 110
        64532 => X"78",  -- 120
        64533 => X"74",  -- 116
        64534 => X"62",  -- 98
        64535 => X"69",  -- 105
        64536 => X"72",  -- 114
        64537 => X"6D",  -- 109
        64538 => X"6F",  -- 111
        64539 => X"6D",  -- 109
        64540 => X"77",  -- 119
        64541 => X"79",  -- 121
        64542 => X"68",  -- 104
        64543 => X"6B",  -- 107
        64544 => X"86",  -- 134
        64545 => X"85",  -- 133
        64546 => X"8A",  -- 138
        64547 => X"87",  -- 135
        64548 => X"7B",  -- 123
        64549 => X"7C",  -- 124
        64550 => X"89",  -- 137
        64551 => X"90",  -- 144
        64552 => X"A6",  -- 166
        64553 => X"A7",  -- 167
        64554 => X"46",  -- 70
        64555 => X"0F",  -- 15
        64556 => X"00",  -- 0
        64557 => X"08",  -- 8
        64558 => X"0F",  -- 15
        64559 => X"09",  -- 9
        64560 => X"23",  -- 35
        64561 => X"48",  -- 72
        64562 => X"6D",  -- 109
        64563 => X"7B",  -- 123
        64564 => X"98",  -- 152
        64565 => X"92",  -- 146
        64566 => X"B2",  -- 178
        64567 => X"BC",  -- 188
        64568 => X"AC",  -- 172
        64569 => X"90",  -- 144
        64570 => X"8D",  -- 141
        64571 => X"97",  -- 151
        64572 => X"A5",  -- 165
        64573 => X"A8",  -- 168
        64574 => X"AE",  -- 174
        64575 => X"AB",  -- 171
        64576 => X"BA",  -- 186
        64577 => X"A9",  -- 169
        64578 => X"A2",  -- 162
        64579 => X"A5",  -- 165
        64580 => X"B4",  -- 180
        64581 => X"AC",  -- 172
        64582 => X"84",  -- 132
        64583 => X"71",  -- 113
        64584 => X"7F",  -- 127
        64585 => X"C2",  -- 194
        64586 => X"B8",  -- 184
        64587 => X"7D",  -- 125
        64588 => X"98",  -- 152
        64589 => X"AA",  -- 170
        64590 => X"B4",  -- 180
        64591 => X"C6",  -- 198
        64592 => X"CC",  -- 204
        64593 => X"D2",  -- 210
        64594 => X"D7",  -- 215
        64595 => X"B7",  -- 183
        64596 => X"74",  -- 116
        64597 => X"49",  -- 73
        64598 => X"45",  -- 69
        64599 => X"47",  -- 71
        64600 => X"3B",  -- 59
        64601 => X"34",  -- 52
        64602 => X"26",  -- 38
        64603 => X"28",  -- 40
        64604 => X"38",  -- 56
        64605 => X"3D",  -- 61
        64606 => X"40",  -- 64
        64607 => X"52",  -- 82
        64608 => X"58",  -- 88
        64609 => X"5B",  -- 91
        64610 => X"59",  -- 89
        64611 => X"51",  -- 81
        64612 => X"46",  -- 70
        64613 => X"41",  -- 65
        64614 => X"46",  -- 70
        64615 => X"4B",  -- 75
        64616 => X"40",  -- 64
        64617 => X"3E",  -- 62
        64618 => X"35",  -- 53
        64619 => X"29",  -- 41
        64620 => X"25",  -- 37
        64621 => X"2B",  -- 43
        64622 => X"37",  -- 55
        64623 => X"3E",  -- 62
        64624 => X"39",  -- 57
        64625 => X"30",  -- 48
        64626 => X"3B",  -- 59
        64627 => X"36",  -- 54
        64628 => X"3E",  -- 62
        64629 => X"38",  -- 56
        64630 => X"3E",  -- 62
        64631 => X"32",  -- 50
        64632 => X"38",  -- 56
        64633 => X"3B",  -- 59
        64634 => X"3A",  -- 58
        64635 => X"39",  -- 57
        64636 => X"3D",  -- 61
        64637 => X"47",  -- 71
        64638 => X"4B",  -- 75
        64639 => X"4B",  -- 75
        64640 => X"77",  -- 119
        64641 => X"74",  -- 116
        64642 => X"6C",  -- 108
        64643 => X"6D",  -- 109
        64644 => X"71",  -- 113
        64645 => X"67",  -- 103
        64646 => X"5C",  -- 92
        64647 => X"60",  -- 96
        64648 => X"72",  -- 114
        64649 => X"70",  -- 112
        64650 => X"70",  -- 112
        64651 => X"74",  -- 116
        64652 => X"74",  -- 116
        64653 => X"6F",  -- 111
        64654 => X"69",  -- 105
        64655 => X"67",  -- 103
        64656 => X"69",  -- 105
        64657 => X"71",  -- 113
        64658 => X"6D",  -- 109
        64659 => X"64",  -- 100
        64660 => X"6D",  -- 109
        64661 => X"5B",  -- 91
        64662 => X"80",  -- 128
        64663 => X"79",  -- 121
        64664 => X"63",  -- 99
        64665 => X"5B",  -- 91
        64666 => X"55",  -- 85
        64667 => X"51",  -- 81
        64668 => X"6B",  -- 107
        64669 => X"69",  -- 105
        64670 => X"6C",  -- 108
        64671 => X"42",  -- 66
        64672 => X"61",  -- 97
        64673 => X"3E",  -- 62
        64674 => X"33",  -- 51
        64675 => X"2C",  -- 44
        64676 => X"32",  -- 50
        64677 => X"23",  -- 35
        64678 => X"5E",  -- 94
        64679 => X"62",  -- 98
        64680 => X"86",  -- 134
        64681 => X"71",  -- 113
        64682 => X"55",  -- 85
        64683 => X"3A",  -- 58
        64684 => X"46",  -- 70
        64685 => X"5A",  -- 90
        64686 => X"38",  -- 56
        64687 => X"3D",  -- 61
        64688 => X"65",  -- 101
        64689 => X"7E",  -- 126
        64690 => X"5F",  -- 95
        64691 => X"83",  -- 131
        64692 => X"39",  -- 57
        64693 => X"6D",  -- 109
        64694 => X"62",  -- 98
        64695 => X"4F",  -- 79
        64696 => X"53",  -- 83
        64697 => X"4C",  -- 76
        64698 => X"4A",  -- 74
        64699 => X"48",  -- 72
        64700 => X"3A",  -- 58
        64701 => X"41",  -- 65
        64702 => X"47",  -- 71
        64703 => X"36",  -- 54
        64704 => X"2D",  -- 45
        64705 => X"3C",  -- 60
        64706 => X"3F",  -- 63
        64707 => X"2B",  -- 43
        64708 => X"1A",  -- 26
        64709 => X"18",  -- 24
        64710 => X"1A",  -- 26
        64711 => X"18",  -- 24
        64712 => X"30",  -- 48
        64713 => X"44",  -- 68
        64714 => X"57",  -- 87
        64715 => X"61",  -- 97
        64716 => X"5F",  -- 95
        64717 => X"72",  -- 114
        64718 => X"6D",  -- 109
        64719 => X"6D",  -- 109
        64720 => X"89",  -- 137
        64721 => X"8C",  -- 140
        64722 => X"82",  -- 130
        64723 => X"5C",  -- 92
        64724 => X"57",  -- 87
        64725 => X"81",  -- 129
        64726 => X"9B",  -- 155
        64727 => X"70",  -- 112
        64728 => X"51",  -- 81
        64729 => X"64",  -- 100
        64730 => X"84",  -- 132
        64731 => X"7A",  -- 122
        64732 => X"73",  -- 115
        64733 => X"6A",  -- 106
        64734 => X"68",  -- 104
        64735 => X"64",  -- 100
        64736 => X"65",  -- 101
        64737 => X"77",  -- 119
        64738 => X"66",  -- 102
        64739 => X"96",  -- 150
        64740 => X"9F",  -- 159
        64741 => X"74",  -- 116
        64742 => X"80",  -- 128
        64743 => X"88",  -- 136
        64744 => X"9F",  -- 159
        64745 => X"9B",  -- 155
        64746 => X"A0",  -- 160
        64747 => X"B7",  -- 183
        64748 => X"A9",  -- 169
        64749 => X"88",  -- 136
        64750 => X"90",  -- 144
        64751 => X"A5",  -- 165
        64752 => X"9E",  -- 158
        64753 => X"7F",  -- 127
        64754 => X"6C",  -- 108
        64755 => X"6C",  -- 108
        64756 => X"69",  -- 105
        64757 => X"63",  -- 99
        64758 => X"63",  -- 99
        64759 => X"45",  -- 69
        64760 => X"47",  -- 71
        64761 => X"5E",  -- 94
        64762 => X"43",  -- 67
        64763 => X"4D",  -- 77
        64764 => X"49",  -- 73
        64765 => X"5E",  -- 94
        64766 => X"57",  -- 87
        64767 => X"3C",  -- 60
        64768 => X"38",  -- 56
        64769 => X"55",  -- 85
        64770 => X"72",  -- 114
        64771 => X"57",  -- 87
        64772 => X"56",  -- 86
        64773 => X"81",  -- 129
        64774 => X"57",  -- 87
        64775 => X"62",  -- 98
        64776 => X"64",  -- 100
        64777 => X"86",  -- 134
        64778 => X"76",  -- 118
        64779 => X"62",  -- 98
        64780 => X"5E",  -- 94
        64781 => X"60",  -- 96
        64782 => X"90",  -- 144
        64783 => X"73",  -- 115
        64784 => X"51",  -- 81
        64785 => X"69",  -- 105
        64786 => X"62",  -- 98
        64787 => X"5C",  -- 92
        64788 => X"95",  -- 149
        64789 => X"59",  -- 89
        64790 => X"46",  -- 70
        64791 => X"43",  -- 67
        64792 => X"31",  -- 49
        64793 => X"16",  -- 22
        64794 => X"14",  -- 20
        64795 => X"0F",  -- 15
        64796 => X"60",  -- 96
        64797 => X"11",  -- 17
        64798 => X"5B",  -- 91
        64799 => X"5A",  -- 90
        64800 => X"5E",  -- 94
        64801 => X"18",  -- 24
        64802 => X"1B",  -- 27
        64803 => X"24",  -- 36
        64804 => X"1D",  -- 29
        64805 => X"2A",  -- 42
        64806 => X"27",  -- 39
        64807 => X"28",  -- 40
        64808 => X"2E",  -- 46
        64809 => X"27",  -- 39
        64810 => X"24",  -- 36
        64811 => X"28",  -- 40
        64812 => X"2D",  -- 45
        64813 => X"2D",  -- 45
        64814 => X"2A",  -- 42
        64815 => X"29",  -- 41
        64816 => X"2A",  -- 42
        64817 => X"2A",  -- 42
        64818 => X"2C",  -- 44
        64819 => X"2F",  -- 47
        64820 => X"31",  -- 49
        64821 => X"2F",  -- 47
        64822 => X"27",  -- 39
        64823 => X"21",  -- 33
        64824 => X"27",  -- 39
        64825 => X"2F",  -- 47
        64826 => X"35",  -- 53
        64827 => X"3B",  -- 59
        64828 => X"3F",  -- 63
        64829 => X"42",  -- 66
        64830 => X"41",  -- 65
        64831 => X"3E",  -- 62
        64832 => X"36",  -- 54
        64833 => X"2E",  -- 46
        64834 => X"2E",  -- 46
        64835 => X"3C",  -- 60
        64836 => X"55",  -- 85
        64837 => X"6F",  -- 111
        64838 => X"83",  -- 131
        64839 => X"8E",  -- 142
        64840 => X"86",  -- 134
        64841 => X"73",  -- 115
        64842 => X"5B",  -- 91
        64843 => X"4D",  -- 77
        64844 => X"4F",  -- 79
        64845 => X"51",  -- 81
        64846 => X"4D",  -- 77
        64847 => X"44",  -- 68
        64848 => X"40",  -- 64
        64849 => X"50",  -- 80
        64850 => X"66",  -- 102
        64851 => X"6B",  -- 107
        64852 => X"73",  -- 115
        64853 => X"72",  -- 114
        64854 => X"63",  -- 99
        64855 => X"67",  -- 103
        64856 => X"71",  -- 113
        64857 => X"71",  -- 113
        64858 => X"71",  -- 113
        64859 => X"67",  -- 103
        64860 => X"6A",  -- 106
        64861 => X"71",  -- 113
        64862 => X"6F",  -- 111
        64863 => X"7E",  -- 126
        64864 => X"91",  -- 145
        64865 => X"90",  -- 144
        64866 => X"8C",  -- 140
        64867 => X"7E",  -- 126
        64868 => X"72",  -- 114
        64869 => X"7F",  -- 127
        64870 => X"95",  -- 149
        64871 => X"9D",  -- 157
        64872 => X"A4",  -- 164
        64873 => X"9E",  -- 158
        64874 => X"37",  -- 55
        64875 => X"00",  -- 0
        64876 => X"07",  -- 7
        64877 => X"12",  -- 18
        64878 => X"0A",  -- 10
        64879 => X"03",  -- 3
        64880 => X"0D",  -- 13
        64881 => X"37",  -- 55
        64882 => X"53",  -- 83
        64883 => X"64",  -- 100
        64884 => X"78",  -- 120
        64885 => X"82",  -- 130
        64886 => X"A0",  -- 160
        64887 => X"AA",  -- 170
        64888 => X"92",  -- 146
        64889 => X"80",  -- 128
        64890 => X"88",  -- 136
        64891 => X"9E",  -- 158
        64892 => X"96",  -- 150
        64893 => X"9C",  -- 156
        64894 => X"A3",  -- 163
        64895 => X"9E",  -- 158
        64896 => X"A8",  -- 168
        64897 => X"AE",  -- 174
        64898 => X"A1",  -- 161
        64899 => X"97",  -- 151
        64900 => X"A4",  -- 164
        64901 => X"89",  -- 137
        64902 => X"68",  -- 104
        64903 => X"85",  -- 133
        64904 => X"8B",  -- 139
        64905 => X"C2",  -- 194
        64906 => X"AE",  -- 174
        64907 => X"6A",  -- 106
        64908 => X"80",  -- 128
        64909 => X"9C",  -- 156
        64910 => X"A9",  -- 169
        64911 => X"AE",  -- 174
        64912 => X"B2",  -- 178
        64913 => X"C0",  -- 192
        64914 => X"C4",  -- 196
        64915 => X"A6",  -- 166
        64916 => X"75",  -- 117
        64917 => X"5C",  -- 92
        64918 => X"59",  -- 89
        64919 => X"57",  -- 87
        64920 => X"56",  -- 86
        64921 => X"4B",  -- 75
        64922 => X"37",  -- 55
        64923 => X"31",  -- 49
        64924 => X"36",  -- 54
        64925 => X"37",  -- 55
        64926 => X"3F",  -- 63
        64927 => X"51",  -- 81
        64928 => X"5A",  -- 90
        64929 => X"59",  -- 89
        64930 => X"50",  -- 80
        64931 => X"42",  -- 66
        64932 => X"3C",  -- 60
        64933 => X"40",  -- 64
        64934 => X"42",  -- 66
        64935 => X"3F",  -- 63
        64936 => X"45",  -- 69
        64937 => X"3A",  -- 58
        64938 => X"2D",  -- 45
        64939 => X"26",  -- 38
        64940 => X"27",  -- 39
        64941 => X"2B",  -- 43
        64942 => X"31",  -- 49
        64943 => X"36",  -- 54
        64944 => X"3D",  -- 61
        64945 => X"34",  -- 52
        64946 => X"3C",  -- 60
        64947 => X"3B",  -- 59
        64948 => X"42",  -- 66
        64949 => X"3E",  -- 62
        64950 => X"41",  -- 65
        64951 => X"34",  -- 52
        64952 => X"27",  -- 39
        64953 => X"2D",  -- 45
        64954 => X"31",  -- 49
        64955 => X"34",  -- 52
        64956 => X"37",  -- 55
        64957 => X"3E",  -- 62
        64958 => X"44",  -- 68
        64959 => X"45",  -- 69
        64960 => X"74",  -- 116
        64961 => X"70",  -- 112
        64962 => X"6C",  -- 108
        64963 => X"6C",  -- 108
        64964 => X"6C",  -- 108
        64965 => X"67",  -- 103
        64966 => X"65",  -- 101
        64967 => X"6A",  -- 106
        64968 => X"73",  -- 115
        64969 => X"6C",  -- 108
        64970 => X"6B",  -- 107
        64971 => X"72",  -- 114
        64972 => X"74",  -- 116
        64973 => X"6D",  -- 109
        64974 => X"66",  -- 102
        64975 => X"65",  -- 101
        64976 => X"6A",  -- 106
        64977 => X"6C",  -- 108
        64978 => X"72",  -- 114
        64979 => X"66",  -- 102
        64980 => X"5B",  -- 91
        64981 => X"73",  -- 115
        64982 => X"8F",  -- 143
        64983 => X"60",  -- 96
        64984 => X"6B",  -- 107
        64985 => X"50",  -- 80
        64986 => X"49",  -- 73
        64987 => X"51",  -- 81
        64988 => X"69",  -- 105
        64989 => X"6A",  -- 106
        64990 => X"65",  -- 101
        64991 => X"48",  -- 72
        64992 => X"6F",  -- 111
        64993 => X"3C",  -- 60
        64994 => X"49",  -- 73
        64995 => X"3C",  -- 60
        64996 => X"3F",  -- 63
        64997 => X"49",  -- 73
        64998 => X"5E",  -- 94
        64999 => X"4E",  -- 78
        65000 => X"66",  -- 102
        65001 => X"4E",  -- 78
        65002 => X"32",  -- 50
        65003 => X"2E",  -- 46
        65004 => X"57",  -- 87
        65005 => X"3A",  -- 58
        65006 => X"3E",  -- 62
        65007 => X"64",  -- 100
        65008 => X"6B",  -- 107
        65009 => X"69",  -- 105
        65010 => X"6A",  -- 106
        65011 => X"4D",  -- 77
        65012 => X"5A",  -- 90
        65013 => X"7F",  -- 127
        65014 => X"40",  -- 64
        65015 => X"4C",  -- 76
        65016 => X"52",  -- 82
        65017 => X"41",  -- 65
        65018 => X"52",  -- 82
        65019 => X"3B",  -- 59
        65020 => X"34",  -- 52
        65021 => X"34",  -- 52
        65022 => X"3A",  -- 58
        65023 => X"3E",  -- 62
        65024 => X"39",  -- 57
        65025 => X"3D",  -- 61
        65026 => X"40",  -- 64
        65027 => X"37",  -- 55
        65028 => X"29",  -- 41
        65029 => X"23",  -- 35
        65030 => X"2D",  -- 45
        65031 => X"3A",  -- 58
        65032 => X"4C",  -- 76
        65033 => X"4E",  -- 78
        65034 => X"54",  -- 84
        65035 => X"4E",  -- 78
        65036 => X"4E",  -- 78
        65037 => X"56",  -- 86
        65038 => X"5B",  -- 91
        65039 => X"75",  -- 117
        65040 => X"92",  -- 146
        65041 => X"94",  -- 148
        65042 => X"66",  -- 102
        65043 => X"55",  -- 85
        65044 => X"89",  -- 137
        65045 => X"8A",  -- 138
        65046 => X"84",  -- 132
        65047 => X"65",  -- 101
        65048 => X"68",  -- 104
        65049 => X"67",  -- 103
        65050 => X"82",  -- 130
        65051 => X"6F",  -- 111
        65052 => X"8B",  -- 139
        65053 => X"80",  -- 128
        65054 => X"6C",  -- 108
        65055 => X"66",  -- 102
        65056 => X"6C",  -- 108
        65057 => X"7E",  -- 126
        65058 => X"86",  -- 134
        65059 => X"87",  -- 135
        65060 => X"9F",  -- 159
        65061 => X"99",  -- 153
        65062 => X"99",  -- 153
        65063 => X"8B",  -- 139
        65064 => X"8D",  -- 141
        65065 => X"91",  -- 145
        65066 => X"9D",  -- 157
        65067 => X"B2",  -- 178
        65068 => X"B5",  -- 181
        65069 => X"A0",  -- 160
        65070 => X"97",  -- 151
        65071 => X"9C",  -- 156
        65072 => X"8F",  -- 143
        65073 => X"8A",  -- 138
        65074 => X"68",  -- 104
        65075 => X"62",  -- 98
        65076 => X"76",  -- 118
        65077 => X"68",  -- 104
        65078 => X"62",  -- 98
        65079 => X"49",  -- 73
        65080 => X"43",  -- 67
        65081 => X"59",  -- 89
        65082 => X"4B",  -- 75
        65083 => X"4B",  -- 75
        65084 => X"48",  -- 72
        65085 => X"4D",  -- 77
        65086 => X"61",  -- 97
        65087 => X"37",  -- 55
        65088 => X"3D",  -- 61
        65089 => X"56",  -- 86
        65090 => X"67",  -- 103
        65091 => X"60",  -- 96
        65092 => X"5D",  -- 93
        65093 => X"78",  -- 120
        65094 => X"53",  -- 83
        65095 => X"5E",  -- 94
        65096 => X"63",  -- 99
        65097 => X"79",  -- 121
        65098 => X"91",  -- 145
        65099 => X"66",  -- 102
        65100 => X"68",  -- 104
        65101 => X"65",  -- 101
        65102 => X"64",  -- 100
        65103 => X"92",  -- 146
        65104 => X"62",  -- 98
        65105 => X"5B",  -- 91
        65106 => X"6C",  -- 108
        65107 => X"50",  -- 80
        65108 => X"55",  -- 85
        65109 => X"84",  -- 132
        65110 => X"3A",  -- 58
        65111 => X"34",  -- 52
        65112 => X"0B",  -- 11
        65113 => X"16",  -- 22
        65114 => X"04",  -- 4
        65115 => X"07",  -- 7
        65116 => X"34",  -- 52
        65117 => X"51",  -- 81
        65118 => X"11",  -- 17
        65119 => X"57",  -- 87
        65120 => X"64",  -- 100
        65121 => X"4F",  -- 79
        65122 => X"0A",  -- 10
        65123 => X"21",  -- 33
        65124 => X"1A",  -- 26
        65125 => X"26",  -- 38
        65126 => X"27",  -- 39
        65127 => X"18",  -- 24
        65128 => X"1F",  -- 31
        65129 => X"23",  -- 35
        65130 => X"2A",  -- 42
        65131 => X"2C",  -- 44
        65132 => X"28",  -- 40
        65133 => X"23",  -- 35
        65134 => X"25",  -- 37
        65135 => X"2B",  -- 43
        65136 => X"2F",  -- 47
        65137 => X"2D",  -- 45
        65138 => X"2C",  -- 44
        65139 => X"2C",  -- 44
        65140 => X"30",  -- 48
        65141 => X"31",  -- 49
        65142 => X"2C",  -- 44
        65143 => X"22",  -- 34
        65144 => X"27",  -- 39
        65145 => X"2E",  -- 46
        65146 => X"37",  -- 55
        65147 => X"3A",  -- 58
        65148 => X"3D",  -- 61
        65149 => X"40",  -- 64
        65150 => X"3D",  -- 61
        65151 => X"37",  -- 55
        65152 => X"31",  -- 49
        65153 => X"2B",  -- 43
        65154 => X"2D",  -- 45
        65155 => X"3A",  -- 58
        65156 => X"4F",  -- 79
        65157 => X"66",  -- 102
        65158 => X"78",  -- 120
        65159 => X"85",  -- 133
        65160 => X"82",  -- 130
        65161 => X"74",  -- 116
        65162 => X"63",  -- 99
        65163 => X"5E",  -- 94
        65164 => X"60",  -- 96
        65165 => X"5F",  -- 95
        65166 => X"53",  -- 83
        65167 => X"48",  -- 72
        65168 => X"41",  -- 65
        65169 => X"4B",  -- 75
        65170 => X"63",  -- 99
        65171 => X"6B",  -- 107
        65172 => X"71",  -- 113
        65173 => X"6B",  -- 107
        65174 => X"59",  -- 89
        65175 => X"5E",  -- 94
        65176 => X"61",  -- 97
        65177 => X"69",  -- 105
        65178 => X"6C",  -- 108
        65179 => X"59",  -- 89
        65180 => X"57",  -- 87
        65181 => X"67",  -- 103
        65182 => X"79",  -- 121
        65183 => X"96",  -- 150
        65184 => X"9B",  -- 155
        65185 => X"95",  -- 149
        65186 => X"8F",  -- 143
        65187 => X"80",  -- 128
        65188 => X"71",  -- 113
        65189 => X"7B",  -- 123
        65190 => X"94",  -- 148
        65191 => X"A1",  -- 161
        65192 => X"9D",  -- 157
        65193 => X"9F",  -- 159
        65194 => X"4A",  -- 74
        65195 => X"13",  -- 19
        65196 => X"1A",  -- 26
        65197 => X"11",  -- 17
        65198 => X"04",  -- 4
        65199 => X"0C",  -- 12
        65200 => X"05",  -- 5
        65201 => X"19",  -- 25
        65202 => X"1F",  -- 31
        65203 => X"3E",  -- 62
        65204 => X"63",  -- 99
        65205 => X"7A",  -- 122
        65206 => X"82",  -- 130
        65207 => X"7B",  -- 123
        65208 => X"58",  -- 88
        65209 => X"53",  -- 83
        65210 => X"65",  -- 101
        65211 => X"7D",  -- 125
        65212 => X"5E",  -- 94
        65213 => X"6B",  -- 107
        65214 => X"7D",  -- 125
        65215 => X"83",  -- 131
        65216 => X"66",  -- 102
        65217 => X"82",  -- 130
        65218 => X"80",  -- 128
        65219 => X"6D",  -- 109
        65220 => X"7B",  -- 123
        65221 => X"79",  -- 121
        65222 => X"6A",  -- 106
        65223 => X"87",  -- 135
        65224 => X"84",  -- 132
        65225 => X"A4",  -- 164
        65226 => X"8B",  -- 139
        65227 => X"4A",  -- 74
        65228 => X"5B",  -- 91
        65229 => X"72",  -- 114
        65230 => X"7F",  -- 127
        65231 => X"7F",  -- 127
        65232 => X"89",  -- 137
        65233 => X"8E",  -- 142
        65234 => X"94",  -- 148
        65235 => X"93",  -- 147
        65236 => X"8E",  -- 142
        65237 => X"8D",  -- 141
        65238 => X"8C",  -- 140
        65239 => X"85",  -- 133
        65240 => X"8E",  -- 142
        65241 => X"8A",  -- 138
        65242 => X"82",  -- 130
        65243 => X"80",  -- 128
        65244 => X"7B",  -- 123
        65245 => X"76",  -- 118
        65246 => X"75",  -- 117
        65247 => X"7B",  -- 123
        65248 => X"78",  -- 120
        65249 => X"78",  -- 120
        65250 => X"72",  -- 114
        65251 => X"67",  -- 103
        65252 => X"64",  -- 100
        65253 => X"66",  -- 102
        65254 => X"64",  -- 100
        65255 => X"5E",  -- 94
        65256 => X"5F",  -- 95
        65257 => X"4C",  -- 76
        65258 => X"3D",  -- 61
        65259 => X"3E",  -- 62
        65260 => X"46",  -- 70
        65261 => X"47",  -- 71
        65262 => X"41",  -- 65
        65263 => X"3B",  -- 59
        65264 => X"42",  -- 66
        65265 => X"38",  -- 56
        65266 => X"3A",  -- 58
        65267 => X"3B",  -- 59
        65268 => X"3C",  -- 60
        65269 => X"39",  -- 57
        65270 => X"35",  -- 53
        65271 => X"26",  -- 38
        65272 => X"32",  -- 50
        65273 => X"39",  -- 57
        65274 => X"3C",  -- 60
        65275 => X"3B",  -- 59
        65276 => X"39",  -- 57
        65277 => X"3A",  -- 58
        65278 => X"3F",  -- 63
        65279 => X"43",  -- 67
        65280 => X"75",  -- 117
        65281 => X"71",  -- 113
        65282 => X"6F",  -- 111
        65283 => X"6D",  -- 109
        65284 => X"67",  -- 103
        65285 => X"69",  -- 105
        65286 => X"71",  -- 113
        65287 => X"78",  -- 120
        65288 => X"75",  -- 117
        65289 => X"6A",  -- 106
        65290 => X"63",  -- 99
        65291 => X"67",  -- 103
        65292 => X"69",  -- 105
        65293 => X"65",  -- 101
        65294 => X"64",  -- 100
        65295 => X"67",  -- 103
        65296 => X"5F",  -- 95
        65297 => X"6A",  -- 106
        65298 => X"5F",  -- 95
        65299 => X"68",  -- 104
        65300 => X"58",  -- 88
        65301 => X"8F",  -- 143
        65302 => X"6F",  -- 111
        65303 => X"5D",  -- 93
        65304 => X"4D",  -- 77
        65305 => X"49",  -- 73
        65306 => X"5F",  -- 95
        65307 => X"64",  -- 100
        65308 => X"5B",  -- 91
        65309 => X"69",  -- 105
        65310 => X"57",  -- 87
        65311 => X"63",  -- 99
        65312 => X"6A",  -- 106
        65313 => X"55",  -- 85
        65314 => X"5C",  -- 92
        65315 => X"4A",  -- 74
        65316 => X"5A",  -- 90
        65317 => X"82",  -- 130
        65318 => X"3A",  -- 58
        65319 => X"71",  -- 113
        65320 => X"42",  -- 66
        65321 => X"63",  -- 99
        65322 => X"26",  -- 38
        65323 => X"27",  -- 39
        65324 => X"63",  -- 99
        65325 => X"30",  -- 48
        65326 => X"3C",  -- 60
        65327 => X"77",  -- 119
        65328 => X"7A",  -- 122
        65329 => X"52",  -- 82
        65330 => X"61",  -- 97
        65331 => X"33",  -- 51
        65332 => X"7C",  -- 124
        65333 => X"62",  -- 98
        65334 => X"3C",  -- 60
        65335 => X"61",  -- 97
        65336 => X"4B",  -- 75
        65337 => X"46",  -- 70
        65338 => X"59",  -- 89
        65339 => X"2A",  -- 42
        65340 => X"27",  -- 39
        65341 => X"37",  -- 55
        65342 => X"40",  -- 64
        65343 => X"3F",  -- 63
        65344 => X"3C",  -- 60
        65345 => X"3F",  -- 63
        65346 => X"41",  -- 65
        65347 => X"3D",  -- 61
        65348 => X"36",  -- 54
        65349 => X"36",  -- 54
        65350 => X"41",  -- 65
        65351 => X"50",  -- 80
        65352 => X"53",  -- 83
        65353 => X"45",  -- 69
        65354 => X"44",  -- 68
        65355 => X"45",  -- 69
        65356 => X"43",  -- 67
        65357 => X"39",  -- 57
        65358 => X"52",  -- 82
        65359 => X"82",  -- 130
        65360 => X"85",  -- 133
        65361 => X"8B",  -- 139
        65362 => X"5B",  -- 91
        65363 => X"62",  -- 98
        65364 => X"8B",  -- 139
        65365 => X"70",  -- 112
        65366 => X"81",  -- 129
        65367 => X"79",  -- 121
        65368 => X"81",  -- 129
        65369 => X"78",  -- 120
        65370 => X"81",  -- 129
        65371 => X"5D",  -- 93
        65372 => X"87",  -- 135
        65373 => X"80",  -- 128
        65374 => X"6B",  -- 107
        65375 => X"5B",  -- 91
        65376 => X"6B",  -- 107
        65377 => X"7D",  -- 125
        65378 => X"91",  -- 145
        65379 => X"89",  -- 137
        65380 => X"99",  -- 153
        65381 => X"9B",  -- 155
        65382 => X"9E",  -- 158
        65383 => X"71",  -- 113
        65384 => X"76",  -- 118
        65385 => X"8D",  -- 141
        65386 => X"9F",  -- 159
        65387 => X"A7",  -- 167
        65388 => X"AF",  -- 175
        65389 => X"A7",  -- 167
        65390 => X"96",  -- 150
        65391 => X"95",  -- 149
        65392 => X"8C",  -- 140
        65393 => X"83",  -- 131
        65394 => X"73",  -- 115
        65395 => X"64",  -- 100
        65396 => X"66",  -- 102
        65397 => X"5F",  -- 95
        65398 => X"6B",  -- 107
        65399 => X"3C",  -- 60
        65400 => X"41",  -- 65
        65401 => X"4E",  -- 78
        65402 => X"54",  -- 84
        65403 => X"47",  -- 71
        65404 => X"4A",  -- 74
        65405 => X"38",  -- 56
        65406 => X"5E",  -- 94
        65407 => X"32",  -- 50
        65408 => X"43",  -- 67
        65409 => X"57",  -- 87
        65410 => X"52",  -- 82
        65411 => X"63",  -- 99
        65412 => X"65",  -- 101
        65413 => X"5F",  -- 95
        65414 => X"4F",  -- 79
        65415 => X"56",  -- 86
        65416 => X"63",  -- 99
        65417 => X"62",  -- 98
        65418 => X"93",  -- 147
        65419 => X"7D",  -- 125
        65420 => X"60",  -- 96
        65421 => X"6D",  -- 109
        65422 => X"50",  -- 80
        65423 => X"7D",  -- 125
        65424 => X"77",  -- 119
        65425 => X"57",  -- 87
        65426 => X"67",  -- 103
        65427 => X"5E",  -- 94
        65428 => X"32",  -- 50
        65429 => X"50",  -- 80
        65430 => X"53",  -- 83
        65431 => X"03",  -- 3
        65432 => X"15",  -- 21
        65433 => X"02",  -- 2
        65434 => X"0A",  -- 10
        65435 => X"0D",  -- 13
        65436 => X"18",  -- 24
        65437 => X"63",  -- 99
        65438 => X"31",  -- 49
        65439 => X"1B",  -- 27
        65440 => X"5A",  -- 90
        65441 => X"76",  -- 118
        65442 => X"2B",  -- 43
        65443 => X"0F",  -- 15
        65444 => X"1F",  -- 31
        65445 => X"1B",  -- 27
        65446 => X"20",  -- 32
        65447 => X"26",  -- 38
        65448 => X"1D",  -- 29
        65449 => X"20",  -- 32
        65450 => X"26",  -- 38
        65451 => X"29",  -- 41
        65452 => X"26",  -- 38
        65453 => X"23",  -- 35
        65454 => X"25",  -- 37
        65455 => X"2B",  -- 43
        65456 => X"2F",  -- 47
        65457 => X"30",  -- 48
        65458 => X"2F",  -- 47
        65459 => X"32",  -- 50
        65460 => X"36",  -- 54
        65461 => X"39",  -- 57
        65462 => X"33",  -- 51
        65463 => X"2A",  -- 42
        65464 => X"25",  -- 37
        65465 => X"2B",  -- 43
        65466 => X"34",  -- 52
        65467 => X"38",  -- 56
        65468 => X"3B",  -- 59
        65469 => X"3C",  -- 60
        65470 => X"3A",  -- 58
        65471 => X"34",  -- 52
        65472 => X"2C",  -- 44
        65473 => X"2C",  -- 44
        65474 => X"31",  -- 49
        65475 => X"3C",  -- 60
        65476 => X"4A",  -- 74
        65477 => X"59",  -- 89
        65478 => X"68",  -- 104
        65479 => X"75",  -- 117
        65480 => X"76",  -- 118
        65481 => X"6C",  -- 108
        65482 => X"63",  -- 99
        65483 => X"65",  -- 101
        65484 => X"6A",  -- 106
        65485 => X"66",  -- 102
        65486 => X"57",  -- 87
        65487 => X"48",  -- 72
        65488 => X"49",  -- 73
        65489 => X"47",  -- 71
        65490 => X"5B",  -- 91
        65491 => X"6A",  -- 106
        65492 => X"6C",  -- 108
        65493 => X"57",  -- 87
        65494 => X"40",  -- 64
        65495 => X"4B",  -- 75
        65496 => X"57",  -- 87
        65497 => X"5C",  -- 92
        65498 => X"5D",  -- 93
        65499 => X"4C",  -- 76
        65500 => X"52",  -- 82
        65501 => X"6B",  -- 107
        65502 => X"7C",  -- 124
        65503 => X"93",  -- 147
        65504 => X"82",  -- 130
        65505 => X"79",  -- 121
        65506 => X"78",  -- 120
        65507 => X"75",  -- 117
        65508 => X"66",  -- 102
        65509 => X"66",  -- 102
        65510 => X"7B",  -- 123
        65511 => X"8E",  -- 142
        65512 => X"97",  -- 151
        65513 => X"A9",  -- 169
        65514 => X"65",  -- 101
        65515 => X"1B",  -- 27
        65516 => X"17",  -- 23
        65517 => X"0F",  -- 15
        65518 => X"09",  -- 9
        65519 => X"17",  -- 23
        65520 => X"0D",  -- 13
        65521 => X"13",  -- 19
        65522 => X"11",  -- 17
        65523 => X"31",  -- 49
        65524 => X"4F",  -- 79
        65525 => X"5C",  -- 92
        65526 => X"63",  -- 99
        65527 => X"67",  -- 103
        65528 => X"4E",  -- 78
        65529 => X"4B",  -- 75
        65530 => X"62",  -- 98
        65531 => X"7B",  -- 123
        65532 => X"5B",  -- 91
        65533 => X"6B",  -- 107
        65534 => X"81",  -- 129
        65535 => X"88",  -- 136
        65536 => X"92",  -- 146
        65537 => X"95",  -- 149
        65538 => X"93",  -- 147
        65539 => X"87",  -- 135
        65540 => X"96",  -- 150
        65541 => X"A8",  -- 168
        65542 => X"9B",  -- 155
        65543 => X"95",  -- 149
        65544 => X"93",  -- 147
        65545 => X"A4",  -- 164
        65546 => X"9B",  -- 155
        65547 => X"7A",  -- 122
        65548 => X"8B",  -- 139
        65549 => X"90",  -- 144
        65550 => X"92",  -- 146
        65551 => X"8C",  -- 140
        65552 => X"8A",  -- 138
        65553 => X"88",  -- 136
        65554 => X"89",  -- 137
        65555 => X"95",  -- 149
        65556 => X"A0",  -- 160
        65557 => X"9F",  -- 159
        65558 => X"99",  -- 153
        65559 => X"98",  -- 152
        65560 => X"85",  -- 133
        65561 => X"8A",  -- 138
        65562 => X"96",  -- 150
        65563 => X"9E",  -- 158
        65564 => X"99",  -- 153
        65565 => X"8F",  -- 143
        65566 => X"89",  -- 137
        65567 => X"83",  -- 131
        65568 => X"86",  -- 134
        65569 => X"8C",  -- 140
        65570 => X"8D",  -- 141
        65571 => X"88",  -- 136
        65572 => X"88",  -- 136
        65573 => X"8F",  -- 143
        65574 => X"90",  -- 144
        65575 => X"8D",  -- 141
        65576 => X"95",  -- 149
        65577 => X"89",  -- 137
        65578 => X"80",  -- 128
        65579 => X"81",  -- 129
        65580 => X"85",  -- 133
        65581 => X"82",  -- 130
        65582 => X"79",  -- 121
        65583 => X"6F",  -- 111
        65584 => X"67",  -- 103
        65585 => X"5D",  -- 93
        65586 => X"59",  -- 89
        65587 => X"5B",  -- 91
        65588 => X"54",  -- 84
        65589 => X"51",  -- 81
        65590 => X"48",  -- 72
        65591 => X"3B",  -- 59
        65592 => X"2D",  -- 45
        65593 => X"31",  -- 49
        65594 => X"35",  -- 53
        65595 => X"36",  -- 54
        65596 => X"34",  -- 52
        65597 => X"36",  -- 54
        65598 => X"3F",  -- 63
        65599 => X"47",  -- 71
        65600 => X"79",  -- 121
        65601 => X"72",  -- 114
        65602 => X"73",  -- 115
        65603 => X"70",  -- 112
        65604 => X"67",  -- 103
        65605 => X"6A",  -- 106
        65606 => X"75",  -- 117
        65607 => X"77",  -- 119
        65608 => X"70",  -- 112
        65609 => X"6E",  -- 110
        65610 => X"6F",  -- 111
        65611 => X"73",  -- 115
        65612 => X"72",  -- 114
        65613 => X"6A",  -- 106
        65614 => X"61",  -- 97
        65615 => X"5C",  -- 92
        65616 => X"4C",  -- 76
        65617 => X"4D",  -- 77
        65618 => X"4F",  -- 79
        65619 => X"46",  -- 70
        65620 => X"77",  -- 119
        65621 => X"6A",  -- 106
        65622 => X"40",  -- 64
        65623 => X"58",  -- 88
        65624 => X"4B",  -- 75
        65625 => X"5D",  -- 93
        65626 => X"70",  -- 112
        65627 => X"5E",  -- 94
        65628 => X"4E",  -- 78
        65629 => X"6D",  -- 109
        65630 => X"58",  -- 88
        65631 => X"76",  -- 118
        65632 => X"64",  -- 100
        65633 => X"5E",  -- 94
        65634 => X"58",  -- 88
        65635 => X"5D",  -- 93
        65636 => X"77",  -- 119
        65637 => X"5B",  -- 91
        65638 => X"68",  -- 104
        65639 => X"83",  -- 131
        65640 => X"50",  -- 80
        65641 => X"59",  -- 89
        65642 => X"1F",  -- 31
        65643 => X"4E",  -- 78
        65644 => X"4E",  -- 78
        65645 => X"31",  -- 49
        65646 => X"41",  -- 65
        65647 => X"70",  -- 112
        65648 => X"6C",  -- 108
        65649 => X"44",  -- 68
        65650 => X"4D",  -- 77
        65651 => X"64",  -- 100
        65652 => X"7C",  -- 124
        65653 => X"34",  -- 52
        65654 => X"4C",  -- 76
        65655 => X"5E",  -- 94
        65656 => X"50",  -- 80
        65657 => X"41",  -- 65
        65658 => X"47",  -- 71
        65659 => X"2A",  -- 42
        65660 => X"33",  -- 51
        65661 => X"3A",  -- 58
        65662 => X"3E",  -- 62
        65663 => X"45",  -- 69
        65664 => X"39",  -- 57
        65665 => X"44",  -- 68
        65666 => X"46",  -- 70
        65667 => X"3B",  -- 59
        65668 => X"3B",  -- 59
        65669 => X"46",  -- 70
        65670 => X"4D",  -- 77
        65671 => X"4A",  -- 74
        65672 => X"48",  -- 72
        65673 => X"3A",  -- 58
        65674 => X"3A",  -- 58
        65675 => X"48",  -- 72
        65676 => X"49",  -- 73
        65677 => X"37",  -- 55
        65678 => X"62",  -- 98
        65679 => X"8A",  -- 138
        65680 => X"6D",  -- 109
        65681 => X"61",  -- 97
        65682 => X"59",  -- 89
        65683 => X"77",  -- 119
        65684 => X"77",  -- 119
        65685 => X"69",  -- 105
        65686 => X"8D",  -- 141
        65687 => X"7B",  -- 123
        65688 => X"83",  -- 131
        65689 => X"89",  -- 137
        65690 => X"86",  -- 134
        65691 => X"53",  -- 83
        65692 => X"71",  -- 113
        65693 => X"77",  -- 119
        65694 => X"74",  -- 116
        65695 => X"5D",  -- 93
        65696 => X"67",  -- 103
        65697 => X"7B",  -- 123
        65698 => X"7D",  -- 125
        65699 => X"8E",  -- 142
        65700 => X"93",  -- 147
        65701 => X"7E",  -- 126
        65702 => X"9F",  -- 159
        65703 => X"78",  -- 120
        65704 => X"6B",  -- 107
        65705 => X"85",  -- 133
        65706 => X"9C",  -- 156
        65707 => X"9E",  -- 158
        65708 => X"A1",  -- 161
        65709 => X"98",  -- 152
        65710 => X"8A",  -- 138
        65711 => X"9C",  -- 156
        65712 => X"7D",  -- 125
        65713 => X"7F",  -- 127
        65714 => X"75",  -- 117
        65715 => X"52",  -- 82
        65716 => X"5E",  -- 94
        65717 => X"5C",  -- 92
        65718 => X"64",  -- 100
        65719 => X"43",  -- 67
        65720 => X"41",  -- 65
        65721 => X"46",  -- 70
        65722 => X"5A",  -- 90
        65723 => X"48",  -- 72
        65724 => X"45",  -- 69
        65725 => X"27",  -- 39
        65726 => X"4A",  -- 74
        65727 => X"36",  -- 54
        65728 => X"47",  -- 71
        65729 => X"53",  -- 83
        65730 => X"48",  -- 72
        65731 => X"5F",  -- 95
        65732 => X"6F",  -- 111
        65733 => X"50",  -- 80
        65734 => X"51",  -- 81
        65735 => X"55",  -- 85
        65736 => X"5D",  -- 93
        65737 => X"57",  -- 87
        65738 => X"7C",  -- 124
        65739 => X"94",  -- 148
        65740 => X"55",  -- 85
        65741 => X"65",  -- 101
        65742 => X"62",  -- 98
        65743 => X"4D",  -- 77
        65744 => X"89",  -- 137
        65745 => X"46",  -- 70
        65746 => X"60",  -- 96
        65747 => X"52",  -- 82
        65748 => X"2D",  -- 45
        65749 => X"0A",  -- 10
        65750 => X"5F",  -- 95
        65751 => X"1A",  -- 26
        65752 => X"0C",  -- 12
        65753 => X"05",  -- 5
        65754 => X"00",  -- 0
        65755 => X"13",  -- 19
        65756 => X"0E",  -- 14
        65757 => X"32",  -- 50
        65758 => X"69",  -- 105
        65759 => X"12",  -- 18
        65760 => X"36",  -- 54
        65761 => X"6F",  -- 111
        65762 => X"76",  -- 118
        65763 => X"01",  -- 1
        65764 => X"0E",  -- 14
        65765 => X"1D",  -- 29
        65766 => X"25",  -- 37
        65767 => X"2E",  -- 46
        65768 => X"2D",  -- 45
        65769 => X"23",  -- 35
        65770 => X"1C",  -- 28
        65771 => X"20",  -- 32
        65772 => X"28",  -- 40
        65773 => X"2C",  -- 44
        65774 => X"2B",  -- 43
        65775 => X"2B",  -- 43
        65776 => X"25",  -- 37
        65777 => X"2A",  -- 42
        65778 => X"2B",  -- 43
        65779 => X"2C",  -- 44
        65780 => X"31",  -- 49
        65781 => X"35",  -- 53
        65782 => X"2F",  -- 47
        65783 => X"26",  -- 38
        65784 => X"24",  -- 36
        65785 => X"2A",  -- 42
        65786 => X"31",  -- 49
        65787 => X"37",  -- 55
        65788 => X"3A",  -- 58
        65789 => X"3F",  -- 63
        65790 => X"3D",  -- 61
        65791 => X"3A",  -- 58
        65792 => X"2D",  -- 45
        65793 => X"31",  -- 49
        65794 => X"38",  -- 56
        65795 => X"42",  -- 66
        65796 => X"49",  -- 73
        65797 => X"51",  -- 81
        65798 => X"5D",  -- 93
        65799 => X"69",  -- 105
        65800 => X"68",  -- 104
        65801 => X"60",  -- 96
        65802 => X"5F",  -- 95
        65803 => X"66",  -- 102
        65804 => X"6E",  -- 110
        65805 => X"69",  -- 105
        65806 => X"59",  -- 89
        65807 => X"4A",  -- 74
        65808 => X"43",  -- 67
        65809 => X"3F",  -- 63
        65810 => X"52",  -- 82
        65811 => X"62",  -- 98
        65812 => X"61",  -- 97
        65813 => X"46",  -- 70
        65814 => X"2F",  -- 47
        65815 => X"43",  -- 67
        65816 => X"5E",  -- 94
        65817 => X"59",  -- 89
        65818 => X"4F",  -- 79
        65819 => X"41",  -- 65
        65820 => X"52",  -- 82
        65821 => X"6C",  -- 108
        65822 => X"68",  -- 104
        65823 => X"67",  -- 103
        65824 => X"58",  -- 88
        65825 => X"56",  -- 86
        65826 => X"62",  -- 98
        65827 => X"6D",  -- 109
        65828 => X"65",  -- 101
        65829 => X"62",  -- 98
        65830 => X"75",  -- 117
        65831 => X"8A",  -- 138
        65832 => X"94",  -- 148
        65833 => X"B6",  -- 182
        65834 => X"89",  -- 137
        65835 => X"2D",  -- 45
        65836 => X"1D",  -- 29
        65837 => X"16",  -- 22
        65838 => X"0A",  -- 10
        65839 => X"06",  -- 6
        65840 => X"05",  -- 5
        65841 => X"15",  -- 21
        65842 => X"22",  -- 34
        65843 => X"34",  -- 52
        65844 => X"47",  -- 71
        65845 => X"47",  -- 71
        65846 => X"69",  -- 105
        65847 => X"83",  -- 131
        65848 => X"8C",  -- 140
        65849 => X"83",  -- 131
        65850 => X"8F",  -- 143
        65851 => X"9D",  -- 157
        65852 => X"8D",  -- 141
        65853 => X"92",  -- 146
        65854 => X"99",  -- 153
        65855 => X"92",  -- 146
        65856 => X"B5",  -- 181
        65857 => X"9F",  -- 159
        65858 => X"A0",  -- 160
        65859 => X"9D",  -- 157
        65860 => X"97",  -- 151
        65861 => X"98",  -- 152
        65862 => X"8E",  -- 142
        65863 => X"8B",  -- 139
        65864 => X"94",  -- 148
        65865 => X"94",  -- 148
        65866 => X"96",  -- 150
        65867 => X"8C",  -- 140
        65868 => X"9B",  -- 155
        65869 => X"96",  -- 150
        65870 => X"96",  -- 150
        65871 => X"8F",  -- 143
        65872 => X"97",  -- 151
        65873 => X"9A",  -- 154
        65874 => X"96",  -- 150
        65875 => X"97",  -- 151
        65876 => X"95",  -- 149
        65877 => X"8A",  -- 138
        65878 => X"85",  -- 133
        65879 => X"90",  -- 144
        65880 => X"8C",  -- 140
        65881 => X"89",  -- 137
        65882 => X"8E",  -- 142
        65883 => X"91",  -- 145
        65884 => X"8A",  -- 138
        65885 => X"8B",  -- 139
        65886 => X"91",  -- 145
        65887 => X"8D",  -- 141
        65888 => X"87",  -- 135
        65889 => X"89",  -- 137
        65890 => X"8B",  -- 139
        65891 => X"8C",  -- 140
        65892 => X"8D",  -- 141
        65893 => X"91",  -- 145
        65894 => X"97",  -- 151
        65895 => X"9C",  -- 156
        65896 => X"9D",  -- 157
        65897 => X"A1",  -- 161
        65898 => X"A0",  -- 160
        65899 => X"97",  -- 151
        65900 => X"8D",  -- 141
        65901 => X"86",  -- 134
        65902 => X"80",  -- 128
        65903 => X"7B",  -- 123
        65904 => X"97",  -- 151
        65905 => X"90",  -- 144
        65906 => X"8C",  -- 140
        65907 => X"94",  -- 148
        65908 => X"8A",  -- 138
        65909 => X"90",  -- 144
        65910 => X"88",  -- 136
        65911 => X"7F",  -- 127
        65912 => X"78",  -- 120
        65913 => X"74",  -- 116
        65914 => X"6C",  -- 108
        65915 => X"60",  -- 96
        65916 => X"51",  -- 81
        65917 => X"45",  -- 69
        65918 => X"44",  -- 68
        65919 => X"48",  -- 72
        65920 => X"74",  -- 116
        65921 => X"6B",  -- 107
        65922 => X"6F",  -- 111
        65923 => X"71",  -- 113
        65924 => X"6B",  -- 107
        65925 => X"70",  -- 112
        65926 => X"75",  -- 117
        65927 => X"6D",  -- 109
        65928 => X"67",  -- 103
        65929 => X"6F",  -- 111
        65930 => X"75",  -- 117
        65931 => X"75",  -- 117
        65932 => X"6E",  -- 110
        65933 => X"63",  -- 99
        65934 => X"53",  -- 83
        65935 => X"46",  -- 70
        65936 => X"3B",  -- 59
        65937 => X"2D",  -- 45
        65938 => X"44",  -- 68
        65939 => X"3F",  -- 63
        65940 => X"6C",  -- 108
        65941 => X"31",  -- 49
        65942 => X"2C",  -- 44
        65943 => X"40",  -- 64
        65944 => X"50",  -- 80
        65945 => X"5D",  -- 93
        65946 => X"56",  -- 86
        65947 => X"47",  -- 71
        65948 => X"59",  -- 89
        65949 => X"6B",  -- 107
        65950 => X"61",  -- 97
        65951 => X"7B",  -- 123
        65952 => X"5F",  -- 95
        65953 => X"55",  -- 85
        65954 => X"53",  -- 83
        65955 => X"6D",  -- 109
        65956 => X"6E",  -- 110
        65957 => X"3C",  -- 60
        65958 => X"90",  -- 144
        65959 => X"6C",  -- 108
        65960 => X"66",  -- 102
        65961 => X"3A",  -- 58
        65962 => X"3D",  -- 61
        65963 => X"79",  -- 121
        65964 => X"47",  -- 71
        65965 => X"50",  -- 80
        65966 => X"73",  -- 115
        65967 => X"87",  -- 135
        65968 => X"50",  -- 80
        65969 => X"53",  -- 83
        65970 => X"55",  -- 85
        65971 => X"8C",  -- 140
        65972 => X"63",  -- 99
        65973 => X"35",  -- 53
        65974 => X"5A",  -- 90
        65975 => X"4A",  -- 74
        65976 => X"53",  -- 83
        65977 => X"45",  -- 69
        65978 => X"42",  -- 66
        65979 => X"3B",  -- 59
        65980 => X"45",  -- 69
        65981 => X"3E",  -- 62
        65982 => X"3F",  -- 63
        65983 => X"4B",  -- 75
        65984 => X"40",  -- 64
        65985 => X"44",  -- 68
        65986 => X"45",  -- 69
        65987 => X"44",  -- 68
        65988 => X"48",  -- 72
        65989 => X"4D",  -- 77
        65990 => X"4A",  -- 74
        65991 => X"41",  -- 65
        65992 => X"40",  -- 64
        65993 => X"44",  -- 68
        65994 => X"3F",  -- 63
        65995 => X"4D",  -- 77
        65996 => X"4E",  -- 78
        65997 => X"41",  -- 65
        65998 => X"79",  -- 121
        65999 => X"7A",  -- 122
        66000 => X"5C",  -- 92
        66001 => X"36",  -- 54
        66002 => X"51",  -- 81
        66003 => X"7E",  -- 126
        66004 => X"75",  -- 117
        66005 => X"79",  -- 121
        66006 => X"7D",  -- 125
        66007 => X"7C",  -- 124
        66008 => X"81",  -- 129
        66009 => X"8B",  -- 139
        66010 => X"7E",  -- 126
        66011 => X"57",  -- 87
        66012 => X"63",  -- 99
        66013 => X"64",  -- 100
        66014 => X"75",  -- 117
        66015 => X"64",  -- 100
        66016 => X"5A",  -- 90
        66017 => X"75",  -- 117
        66018 => X"7A",  -- 122
        66019 => X"8A",  -- 138
        66020 => X"8C",  -- 140
        66021 => X"71",  -- 113
        66022 => X"88",  -- 136
        66023 => X"90",  -- 144
        66024 => X"74",  -- 116
        66025 => X"73",  -- 115
        66026 => X"86",  -- 134
        66027 => X"98",  -- 152
        66028 => X"9E",  -- 158
        66029 => X"80",  -- 128
        66030 => X"6B",  -- 107
        66031 => X"95",  -- 149
        66032 => X"78",  -- 120
        66033 => X"70",  -- 112
        66034 => X"76",  -- 118
        66035 => X"4E",  -- 78
        66036 => X"5B",  -- 91
        66037 => X"5A",  -- 90
        66038 => X"5D",  -- 93
        66039 => X"47",  -- 71
        66040 => X"41",  -- 65
        66041 => X"44",  -- 68
        66042 => X"55",  -- 85
        66043 => X"50",  -- 80
        66044 => X"3D",  -- 61
        66045 => X"25",  -- 37
        66046 => X"38",  -- 56
        66047 => X"47",  -- 71
        66048 => X"47",  -- 71
        66049 => X"47",  -- 71
        66050 => X"4C",  -- 76
        66051 => X"55",  -- 85
        66052 => X"74",  -- 116
        66053 => X"56",  -- 86
        66054 => X"58",  -- 88
        66055 => X"5D",  -- 93
        66056 => X"5E",  -- 94
        66057 => X"61",  -- 97
        66058 => X"65",  -- 101
        66059 => X"92",  -- 146
        66060 => X"66",  -- 102
        66061 => X"57",  -- 87
        66062 => X"59",  -- 89
        66063 => X"3E",  -- 62
        66064 => X"6D",  -- 109
        66065 => X"50",  -- 80
        66066 => X"32",  -- 50
        66067 => X"55",  -- 85
        66068 => X"0B",  -- 11
        66069 => X"0D",  -- 13
        66070 => X"27",  -- 39
        66071 => X"63",  -- 99
        66072 => X"10",  -- 16
        66073 => X"07",  -- 7
        66074 => X"04",  -- 4
        66075 => X"00",  -- 0
        66076 => X"15",  -- 21
        66077 => X"05",  -- 5
        66078 => X"5A",  -- 90
        66079 => X"43",  -- 67
        66080 => X"1B",  -- 27
        66081 => X"3D",  -- 61
        66082 => X"83",  -- 131
        66083 => X"34",  -- 52
        66084 => X"06",  -- 6
        66085 => X"1D",  -- 29
        66086 => X"2A",  -- 42
        66087 => X"27",  -- 39
        66088 => X"31",  -- 49
        66089 => X"24",  -- 36
        66090 => X"1B",  -- 27
        66091 => X"1F",  -- 31
        66092 => X"29",  -- 41
        66093 => X"30",  -- 48
        66094 => X"2E",  -- 46
        66095 => X"2A",  -- 42
        66096 => X"25",  -- 37
        66097 => X"27",  -- 39
        66098 => X"25",  -- 37
        66099 => X"20",  -- 32
        66100 => X"22",  -- 34
        66101 => X"29",  -- 41
        66102 => X"2C",  -- 44
        66103 => X"27",  -- 39
        66104 => X"2D",  -- 45
        66105 => X"32",  -- 50
        66106 => X"36",  -- 54
        66107 => X"39",  -- 57
        66108 => X"3D",  -- 61
        66109 => X"40",  -- 64
        66110 => X"41",  -- 65
        66111 => X"3D",  -- 61
        66112 => X"38",  -- 56
        66113 => X"39",  -- 57
        66114 => X"3E",  -- 62
        66115 => X"47",  -- 71
        66116 => X"4E",  -- 78
        66117 => X"54",  -- 84
        66118 => X"5D",  -- 93
        66119 => X"64",  -- 100
        66120 => X"63",  -- 99
        66121 => X"5B",  -- 91
        66122 => X"5A",  -- 90
        66123 => X"65",  -- 101
        66124 => X"6E",  -- 110
        66125 => X"67",  -- 103
        66126 => X"56",  -- 86
        66127 => X"48",  -- 72
        66128 => X"3D",  -- 61
        66129 => X"41",  -- 65
        66130 => X"54",  -- 84
        66131 => X"5A",  -- 90
        66132 => X"52",  -- 82
        66133 => X"3B",  -- 59
        66134 => X"2E",  -- 46
        66135 => X"44",  -- 68
        66136 => X"5E",  -- 94
        66137 => X"55",  -- 85
        66138 => X"44",  -- 68
        66139 => X"31",  -- 49
        66140 => X"42",  -- 66
        66141 => X"58",  -- 88
        66142 => X"4C",  -- 76
        66143 => X"42",  -- 66
        66144 => X"46",  -- 70
        66145 => X"4E",  -- 78
        66146 => X"64",  -- 100
        66147 => X"71",  -- 113
        66148 => X"6D",  -- 109
        66149 => X"72",  -- 114
        66150 => X"85",  -- 133
        66151 => X"93",  -- 147
        66152 => X"96",  -- 150
        66153 => X"B7",  -- 183
        66154 => X"A8",  -- 168
        66155 => X"5A",  -- 90
        66156 => X"3B",  -- 59
        66157 => X"1E",  -- 30
        66158 => X"10",  -- 16
        66159 => X"0E",  -- 14
        66160 => X"20",  -- 32
        66161 => X"2B",  -- 43
        66162 => X"3A",  -- 58
        66163 => X"47",  -- 71
        66164 => X"6E",  -- 110
        66165 => X"72",  -- 114
        66166 => X"90",  -- 144
        66167 => X"97",  -- 151
        66168 => X"A1",  -- 161
        66169 => X"93",  -- 147
        66170 => X"97",  -- 151
        66171 => X"97",  -- 151
        66172 => X"96",  -- 150
        66173 => X"8F",  -- 143
        66174 => X"91",  -- 145
        66175 => X"86",  -- 134
        66176 => X"98",  -- 152
        66177 => X"8B",  -- 139
        66178 => X"94",  -- 148
        66179 => X"96",  -- 150
        66180 => X"8C",  -- 140
        66181 => X"84",  -- 132
        66182 => X"85",  -- 133
        66183 => X"9A",  -- 154
        66184 => X"9C",  -- 156
        66185 => X"8F",  -- 143
        66186 => X"8E",  -- 142
        66187 => X"86",  -- 134
        66188 => X"91",  -- 145
        66189 => X"8D",  -- 141
        66190 => X"93",  -- 147
        66191 => X"8C",  -- 140
        66192 => X"81",  -- 129
        66193 => X"91",  -- 145
        66194 => X"90",  -- 144
        66195 => X"86",  -- 134
        66196 => X"84",  -- 132
        66197 => X"83",  -- 131
        66198 => X"89",  -- 137
        66199 => X"9C",  -- 156
        66200 => X"97",  -- 151
        66201 => X"8A",  -- 138
        66202 => X"85",  -- 133
        66203 => X"82",  -- 130
        66204 => X"7B",  -- 123
        66205 => X"86",  -- 134
        66206 => X"94",  -- 148
        66207 => X"93",  -- 147
        66208 => X"96",  -- 150
        66209 => X"90",  -- 144
        66210 => X"90",  -- 144
        66211 => X"96",  -- 150
        66212 => X"98",  -- 152
        66213 => X"96",  -- 150
        66214 => X"9A",  -- 154
        66215 => X"A1",  -- 161
        66216 => X"B1",  -- 177
        66217 => X"B5",  -- 181
        66218 => X"B0",  -- 176
        66219 => X"A3",  -- 163
        66220 => X"9C",  -- 156
        66221 => X"9E",  -- 158
        66222 => X"9B",  -- 155
        66223 => X"94",  -- 148
        66224 => X"98",  -- 152
        66225 => X"97",  -- 151
        66226 => X"94",  -- 148
        66227 => X"A2",  -- 162
        66228 => X"98",  -- 152
        66229 => X"A5",  -- 165
        66230 => X"A2",  -- 162
        66231 => X"A1",  -- 161
        66232 => X"A1",  -- 161
        66233 => X"9F",  -- 159
        66234 => X"A0",  -- 160
        66235 => X"9F",  -- 159
        66236 => X"9E",  -- 158
        66237 => X"9D",  -- 157
        66238 => X"A2",  -- 162
        66239 => X"AA",  -- 170
        66240 => X"6A",  -- 106
        66241 => X"60",  -- 96
        66242 => X"67",  -- 103
        66243 => X"71",  -- 113
        66244 => X"71",  -- 113
        66245 => X"77",  -- 119
        66246 => X"77",  -- 119
        66247 => X"65",  -- 101
        66248 => X"64",  -- 100
        66249 => X"68",  -- 104
        66250 => X"64",  -- 100
        66251 => X"56",  -- 86
        66252 => X"4B",  -- 75
        66253 => X"47",  -- 71
        66254 => X"40",  -- 64
        66255 => X"37",  -- 55
        66256 => X"34",  -- 52
        66257 => X"2B",  -- 43
        66258 => X"33",  -- 51
        66259 => X"6C",  -- 108
        66260 => X"31",  -- 49
        66261 => X"24",  -- 36
        66262 => X"2D",  -- 45
        66263 => X"27",  -- 39
        66264 => X"31",  -- 49
        66265 => X"3C",  -- 60
        66266 => X"34",  -- 52
        66267 => X"3F",  -- 63
        66268 => X"6F",  -- 111
        66269 => X"5B",  -- 91
        66270 => X"62",  -- 98
        66271 => X"7F",  -- 127
        66272 => X"55",  -- 85
        66273 => X"54",  -- 84
        66274 => X"59",  -- 89
        66275 => X"70",  -- 112
        66276 => X"48",  -- 72
        66277 => X"74",  -- 116
        66278 => X"5B",  -- 91
        66279 => X"61",  -- 97
        66280 => X"6D",  -- 109
        66281 => X"54",  -- 84
        66282 => X"75",  -- 117
        66283 => X"69",  -- 105
        66284 => X"45",  -- 69
        66285 => X"5F",  -- 95
        66286 => X"7A",  -- 122
        66287 => X"7E",  -- 126
        66288 => X"4B",  -- 75
        66289 => X"73",  -- 115
        66290 => X"71",  -- 113
        66291 => X"84",  -- 132
        66292 => X"4A",  -- 74
        66293 => X"58",  -- 88
        66294 => X"65",  -- 101
        66295 => X"47",  -- 71
        66296 => X"45",  -- 69
        66297 => X"5D",  -- 93
        66298 => X"5A",  -- 90
        66299 => X"43",  -- 67
        66300 => X"43",  -- 67
        66301 => X"4C",  -- 76
        66302 => X"4E",  -- 78
        66303 => X"45",  -- 69
        66304 => X"4B",  -- 75
        66305 => X"3C",  -- 60
        66306 => X"3D",  -- 61
        66307 => X"4F",  -- 79
        66308 => X"56",  -- 86
        66309 => X"48",  -- 72
        66310 => X"3D",  -- 61
        66311 => X"3F",  -- 63
        66312 => X"40",  -- 64
        66313 => X"51",  -- 81
        66314 => X"45",  -- 69
        66315 => X"47",  -- 71
        66316 => X"45",  -- 69
        66317 => X"42",  -- 66
        66318 => X"82",  -- 130
        66319 => X"5F",  -- 95
        66320 => X"55",  -- 85
        66321 => X"28",  -- 40
        66322 => X"4B",  -- 75
        66323 => X"73",  -- 115
        66324 => X"76",  -- 118
        66325 => X"7A",  -- 122
        66326 => X"5B",  -- 91
        66327 => X"98",  -- 152
        66328 => X"8B",  -- 139
        66329 => X"85",  -- 133
        66330 => X"6D",  -- 109
        66331 => X"5E",  -- 94
        66332 => X"5F",  -- 95
        66333 => X"4D",  -- 77
        66334 => X"64",  -- 100
        66335 => X"5E",  -- 94
        66336 => X"46",  -- 70
        66337 => X"6A",  -- 106
        66338 => X"92",  -- 146
        66339 => X"86",  -- 134
        66340 => X"89",  -- 137
        66341 => X"7A",  -- 122
        66342 => X"5C",  -- 92
        66343 => X"8E",  -- 142
        66344 => X"88",  -- 136
        66345 => X"65",  -- 101
        66346 => X"6D",  -- 109
        66347 => X"94",  -- 148
        66348 => X"A4",  -- 164
        66349 => X"70",  -- 112
        66350 => X"49",  -- 73
        66351 => X"7A",  -- 122
        66352 => X"8F",  -- 143
        66353 => X"4F",  -- 79
        66354 => X"80",  -- 128
        66355 => X"6C",  -- 108
        66356 => X"49",  -- 73
        66357 => X"51",  -- 81
        66358 => X"6B",  -- 107
        66359 => X"31",  -- 49
        66360 => X"40",  -- 64
        66361 => X"43",  -- 67
        66362 => X"4F",  -- 79
        66363 => X"58",  -- 88
        66364 => X"37",  -- 55
        66365 => X"2C",  -- 44
        66366 => X"30",  -- 48
        66367 => X"5B",  -- 91
        66368 => X"40",  -- 64
        66369 => X"3A",  -- 58
        66370 => X"52",  -- 82
        66371 => X"4A",  -- 74
        66372 => X"73",  -- 115
        66373 => X"5F",  -- 95
        66374 => X"5A",  -- 90
        66375 => X"61",  -- 97
        66376 => X"65",  -- 101
        66377 => X"70",  -- 112
        66378 => X"5C",  -- 92
        66379 => X"81",  -- 129
        66380 => X"85",  -- 133
        66381 => X"50",  -- 80
        66382 => X"32",  -- 50
        66383 => X"4D",  -- 77
        66384 => X"38",  -- 56
        66385 => X"63",  -- 99
        66386 => X"15",  -- 21
        66387 => X"49",  -- 73
        66388 => X"12",  -- 18
        66389 => X"01",  -- 1
        66390 => X"00",  -- 0
        66391 => X"7A",  -- 122
        66392 => X"3F",  -- 63
        66393 => X"00",  -- 0
        66394 => X"0D",  -- 13
        66395 => X"06",  -- 6
        66396 => X"05",  -- 5
        66397 => X"15",  -- 21
        66398 => X"25",  -- 37
        66399 => X"63",  -- 99
        66400 => X"20",  -- 32
        66401 => X"05",  -- 5
        66402 => X"50",  -- 80
        66403 => X"8F",  -- 143
        66404 => X"1C",  -- 28
        66405 => X"0D",  -- 13
        66406 => X"23",  -- 35
        66407 => X"27",  -- 39
        66408 => X"25",  -- 37
        66409 => X"22",  -- 34
        66410 => X"21",  -- 33
        66411 => X"25",  -- 37
        66412 => X"29",  -- 41
        66413 => X"29",  -- 41
        66414 => X"29",  -- 41
        66415 => X"28",  -- 40
        66416 => X"34",  -- 52
        66417 => X"33",  -- 51
        66418 => X"28",  -- 40
        66419 => X"1B",  -- 27
        66420 => X"1A",  -- 26
        66421 => X"28",  -- 40
        66422 => X"32",  -- 50
        66423 => X"34",  -- 52
        66424 => X"39",  -- 57
        66425 => X"3C",  -- 60
        66426 => X"3E",  -- 62
        66427 => X"3E",  -- 62
        66428 => X"3F",  -- 63
        66429 => X"42",  -- 66
        66430 => X"42",  -- 66
        66431 => X"3F",  -- 63
        66432 => X"42",  -- 66
        66433 => X"3F",  -- 63
        66434 => X"42",  -- 66
        66435 => X"4B",  -- 75
        66436 => X"53",  -- 83
        66437 => X"5B",  -- 91
        66438 => X"60",  -- 96
        66439 => X"66",  -- 102
        66440 => X"63",  -- 99
        66441 => X"5B",  -- 91
        66442 => X"59",  -- 89
        66443 => X"64",  -- 100
        66444 => X"6C",  -- 108
        66445 => X"65",  -- 101
        66446 => X"53",  -- 83
        66447 => X"44",  -- 68
        66448 => X"42",  -- 66
        66449 => X"4D",  -- 77
        66450 => X"5F",  -- 95
        66451 => X"57",  -- 87
        66452 => X"46",  -- 70
        66453 => X"34",  -- 52
        66454 => X"2C",  -- 44
        66455 => X"42",  -- 66
        66456 => X"4A",  -- 74
        66457 => X"45",  -- 69
        66458 => X"38",  -- 56
        66459 => X"1F",  -- 31
        66460 => X"2A",  -- 42
        66461 => X"43",  -- 67
        66462 => X"40",  -- 64
        66463 => X"3F",  -- 63
        66464 => X"4F",  -- 79
        66465 => X"5E",  -- 94
        66466 => X"74",  -- 116
        66467 => X"78",  -- 120
        66468 => X"73",  -- 115
        66469 => X"79",  -- 121
        66470 => X"89",  -- 137
        66471 => X"8E",  -- 142
        66472 => X"9D",  -- 157
        66473 => X"AF",  -- 175
        66474 => X"B6",  -- 182
        66475 => X"82",  -- 130
        66476 => X"59",  -- 89
        66477 => X"24",  -- 36
        66478 => X"21",  -- 33
        66479 => X"3C",  -- 60
        66480 => X"5D",  -- 93
        66481 => X"7C",  -- 124
        66482 => X"94",  -- 148
        66483 => X"82",  -- 130
        66484 => X"8A",  -- 138
        66485 => X"72",  -- 114
        66486 => X"8C",  -- 140
        66487 => X"8C",  -- 140
        66488 => X"91",  -- 145
        66489 => X"8A",  -- 138
        66490 => X"91",  -- 145
        66491 => X"8A",  -- 138
        66492 => X"95",  -- 149
        66493 => X"8D",  -- 141
        66494 => X"99",  -- 153
        66495 => X"9A",  -- 154
        66496 => X"8E",  -- 142
        66497 => X"89",  -- 137
        66498 => X"87",  -- 135
        66499 => X"83",  -- 131
        66500 => X"8B",  -- 139
        66501 => X"89",  -- 137
        66502 => X"81",  -- 129
        66503 => X"96",  -- 150
        66504 => X"A0",  -- 160
        66505 => X"91",  -- 145
        66506 => X"93",  -- 147
        66507 => X"8B",  -- 139
        66508 => X"94",  -- 148
        66509 => X"92",  -- 146
        66510 => X"99",  -- 153
        66511 => X"8C",  -- 140
        66512 => X"84",  -- 132
        66513 => X"98",  -- 152
        66514 => X"91",  -- 145
        66515 => X"7A",  -- 122
        66516 => X"7A",  -- 122
        66517 => X"82",  -- 130
        66518 => X"89",  -- 137
        66519 => X"95",  -- 149
        66520 => X"91",  -- 145
        66521 => X"8A",  -- 138
        66522 => X"92",  -- 146
        66523 => X"99",  -- 153
        66524 => X"94",  -- 148
        66525 => X"9C",  -- 156
        66526 => X"A1",  -- 161
        66527 => X"98",  -- 152
        66528 => X"98",  -- 152
        66529 => X"8E",  -- 142
        66530 => X"91",  -- 145
        66531 => X"9D",  -- 157
        66532 => X"A2",  -- 162
        66533 => X"9A",  -- 154
        66534 => X"99",  -- 153
        66535 => X"9F",  -- 159
        66536 => X"AB",  -- 171
        66537 => X"A9",  -- 169
        66538 => X"9E",  -- 158
        66539 => X"94",  -- 148
        66540 => X"9F",  -- 159
        66541 => X"B2",  -- 178
        66542 => X"B1",  -- 177
        66543 => X"A0",  -- 160
        66544 => X"89",  -- 137
        66545 => X"8A",  -- 138
        66546 => X"86",  -- 134
        66547 => X"95",  -- 149
        66548 => X"88",  -- 136
        66549 => X"97",  -- 151
        66550 => X"96",  -- 150
        66551 => X"96",  -- 150
        66552 => X"A6",  -- 166
        66553 => X"A2",  -- 162
        66554 => X"A3",  -- 163
        66555 => X"A4",  -- 164
        66556 => X"A4",  -- 164
        66557 => X"A1",  -- 161
        66558 => X"A5",  -- 165
        66559 => X"AC",  -- 172
        66560 => X"67",  -- 103
        66561 => X"72",  -- 114
        66562 => X"6D",  -- 109
        66563 => X"6A",  -- 106
        66564 => X"7A",  -- 122
        66565 => X"7A",  -- 122
        66566 => X"6A",  -- 106
        66567 => X"64",  -- 100
        66568 => X"5A",  -- 90
        66569 => X"4E",  -- 78
        66570 => X"3B",  -- 59
        66571 => X"35",  -- 53
        66572 => X"40",  -- 64
        66573 => X"43",  -- 67
        66574 => X"40",  -- 64
        66575 => X"40",  -- 64
        66576 => X"46",  -- 70
        66577 => X"37",  -- 55
        66578 => X"59",  -- 89
        66579 => X"48",  -- 72
        66580 => X"1E",  -- 30
        66581 => X"2F",  -- 47
        66582 => X"38",  -- 56
        66583 => X"28",  -- 40
        66584 => X"21",  -- 33
        66585 => X"38",  -- 56
        66586 => X"47",  -- 71
        66587 => X"62",  -- 98
        66588 => X"78",  -- 120
        66589 => X"58",  -- 88
        66590 => X"6A",  -- 106
        66591 => X"78",  -- 120
        66592 => X"55",  -- 85
        66593 => X"4E",  -- 78
        66594 => X"65",  -- 101
        66595 => X"4D",  -- 77
        66596 => X"59",  -- 89
        66597 => X"87",  -- 135
        66598 => X"51",  -- 81
        66599 => X"7F",  -- 127
        66600 => X"71",  -- 113
        66601 => X"4C",  -- 76
        66602 => X"61",  -- 97
        66603 => X"62",  -- 98
        66604 => X"42",  -- 66
        66605 => X"6F",  -- 111
        66606 => X"92",  -- 146
        66607 => X"53",  -- 83
        66608 => X"60",  -- 96
        66609 => X"6C",  -- 108
        66610 => X"8B",  -- 139
        66611 => X"60",  -- 96
        66612 => X"45",  -- 69
        66613 => X"72",  -- 114
        66614 => X"50",  -- 80
        66615 => X"53",  -- 83
        66616 => X"4E",  -- 78
        66617 => X"69",  -- 105
        66618 => X"52",  -- 82
        66619 => X"4A",  -- 74
        66620 => X"53",  -- 83
        66621 => X"46",  -- 70
        66622 => X"44",  -- 68
        66623 => X"43",  -- 67
        66624 => X"45",  -- 69
        66625 => X"47",  -- 71
        66626 => X"4C",  -- 76
        66627 => X"52",  -- 82
        66628 => X"53",  -- 83
        66629 => X"4B",  -- 75
        66630 => X"42",  -- 66
        66631 => X"3F",  -- 63
        66632 => X"48",  -- 72
        66633 => X"53",  -- 83
        66634 => X"42",  -- 66
        66635 => X"35",  -- 53
        66636 => X"3D",  -- 61
        66637 => X"3E",  -- 62
        66638 => X"68",  -- 104
        66639 => X"4E",  -- 78
        66640 => X"3A",  -- 58
        66641 => X"30",  -- 48
        66642 => X"58",  -- 88
        66643 => X"6C",  -- 108
        66644 => X"72",  -- 114
        66645 => X"64",  -- 100
        66646 => X"4E",  -- 78
        66647 => X"8B",  -- 139
        66648 => X"8D",  -- 141
        66649 => X"6B",  -- 107
        66650 => X"64",  -- 100
        66651 => X"50",  -- 80
        66652 => X"31",  -- 49
        66653 => X"3F",  -- 63
        66654 => X"53",  -- 83
        66655 => X"58",  -- 88
        66656 => X"42",  -- 66
        66657 => X"46",  -- 70
        66658 => X"89",  -- 137
        66659 => X"83",  -- 131
        66660 => X"7E",  -- 126
        66661 => X"6C",  -- 108
        66662 => X"38",  -- 56
        66663 => X"73",  -- 115
        66664 => X"86",  -- 134
        66665 => X"78",  -- 120
        66666 => X"3A",  -- 58
        66667 => X"83",  -- 131
        66668 => X"91",  -- 145
        66669 => X"7B",  -- 123
        66670 => X"3F",  -- 63
        66671 => X"56",  -- 86
        66672 => X"7C",  -- 124
        66673 => X"5B",  -- 91
        66674 => X"68",  -- 104
        66675 => X"71",  -- 113
        66676 => X"53",  -- 83
        66677 => X"50",  -- 80
        66678 => X"57",  -- 87
        66679 => X"3A",  -- 58
        66680 => X"3F",  -- 63
        66681 => X"3B",  -- 59
        66682 => X"42",  -- 66
        66683 => X"4D",  -- 77
        66684 => X"4A",  -- 74
        66685 => X"39",  -- 57
        66686 => X"31",  -- 49
        66687 => X"36",  -- 54
        66688 => X"2B",  -- 43
        66689 => X"37",  -- 55
        66690 => X"45",  -- 69
        66691 => X"54",  -- 84
        66692 => X"72",  -- 114
        66693 => X"5C",  -- 92
        66694 => X"62",  -- 98
        66695 => X"68",  -- 104
        66696 => X"64",  -- 100
        66697 => X"67",  -- 103
        66698 => X"6B",  -- 107
        66699 => X"63",  -- 99
        66700 => X"70",  -- 112
        66701 => X"50",  -- 80
        66702 => X"38",  -- 56
        66703 => X"26",  -- 38
        66704 => X"1C",  -- 28
        66705 => X"43",  -- 67
        66706 => X"0C",  -- 12
        66707 => X"26",  -- 38
        66708 => X"1E",  -- 30
        66709 => X"00",  -- 0
        66710 => X"0F",  -- 15
        66711 => X"16",  -- 22
        66712 => X"7C",  -- 124
        66713 => X"30",  -- 48
        66714 => X"05",  -- 5
        66715 => X"08",  -- 8
        66716 => X"15",  -- 21
        66717 => X"14",  -- 20
        66718 => X"1A",  -- 26
        66719 => X"3D",  -- 61
        66720 => X"53",  -- 83
        66721 => X"11",  -- 17
        66722 => X"17",  -- 23
        66723 => X"73",  -- 115
        66724 => X"41",  -- 65
        66725 => X"0D",  -- 13
        66726 => X"21",  -- 33
        66727 => X"1A",  -- 26
        66728 => X"1D",  -- 29
        66729 => X"26",  -- 38
        66730 => X"2F",  -- 47
        66731 => X"31",  -- 49
        66732 => X"2E",  -- 46
        66733 => X"2B",  -- 43
        66734 => X"2E",  -- 46
        66735 => X"33",  -- 51
        66736 => X"39",  -- 57
        66737 => X"37",  -- 55
        66738 => X"2A",  -- 42
        66739 => X"27",  -- 39
        66740 => X"30",  -- 48
        66741 => X"35",  -- 53
        66742 => X"36",  -- 54
        66743 => X"3C",  -- 60
        66744 => X"40",  -- 64
        66745 => X"3F",  -- 63
        66746 => X"3C",  -- 60
        66747 => X"3E",  -- 62
        66748 => X"46",  -- 70
        66749 => X"4A",  -- 74
        66750 => X"47",  -- 71
        66751 => X"3E",  -- 62
        66752 => X"41",  -- 65
        66753 => X"43",  -- 67
        66754 => X"49",  -- 73
        66755 => X"51",  -- 81
        66756 => X"57",  -- 87
        66757 => X"5C",  -- 92
        66758 => X"65",  -- 101
        66759 => X"6C",  -- 108
        66760 => X"6E",  -- 110
        66761 => X"70",  -- 112
        66762 => X"63",  -- 99
        66763 => X"62",  -- 98
        66764 => X"69",  -- 105
        66765 => X"5B",  -- 91
        66766 => X"43",  -- 67
        66767 => X"3F",  -- 63
        66768 => X"4A",  -- 74
        66769 => X"56",  -- 86
        66770 => X"57",  -- 87
        66771 => X"4A",  -- 74
        66772 => X"3D",  -- 61
        66773 => X"38",  -- 56
        66774 => X"35",  -- 53
        66775 => X"31",  -- 49
        66776 => X"3D",  -- 61
        66777 => X"32",  -- 50
        66778 => X"1F",  -- 31
        66779 => X"11",  -- 17
        66780 => X"14",  -- 20
        66781 => X"25",  -- 37
        66782 => X"34",  -- 52
        66783 => X"3B",  -- 59
        66784 => X"56",  -- 86
        66785 => X"65",  -- 101
        66786 => X"6D",  -- 109
        66787 => X"70",  -- 112
        66788 => X"7E",  -- 126
        66789 => X"77",  -- 119
        66790 => X"6D",  -- 109
        66791 => X"85",  -- 133
        66792 => X"90",  -- 144
        66793 => X"AC",  -- 172
        66794 => X"B8",  -- 184
        66795 => X"9B",  -- 155
        66796 => X"68",  -- 104
        66797 => X"55",  -- 85
        66798 => X"6D",  -- 109
        66799 => X"90",  -- 144
        66800 => X"92",  -- 146
        66801 => X"A0",  -- 160
        66802 => X"8F",  -- 143
        66803 => X"8E",  -- 142
        66804 => X"89",  -- 137
        66805 => X"7C",  -- 124
        66806 => X"89",  -- 137
        66807 => X"8A",  -- 138
        66808 => X"92",  -- 146
        66809 => X"8C",  -- 140
        66810 => X"91",  -- 145
        66811 => X"95",  -- 149
        66812 => X"90",  -- 144
        66813 => X"8E",  -- 142
        66814 => X"90",  -- 144
        66815 => X"8F",  -- 143
        66816 => X"8C",  -- 140
        66817 => X"85",  -- 133
        66818 => X"8C",  -- 140
        66819 => X"91",  -- 145
        66820 => X"8A",  -- 138
        66821 => X"90",  -- 144
        66822 => X"98",  -- 152
        66823 => X"92",  -- 146
        66824 => X"99",  -- 153
        66825 => X"8E",  -- 142
        66826 => X"91",  -- 145
        66827 => X"8D",  -- 141
        66828 => X"9B",  -- 155
        66829 => X"93",  -- 147
        66830 => X"9C",  -- 156
        66831 => X"9B",  -- 155
        66832 => X"97",  -- 151
        66833 => X"91",  -- 145
        66834 => X"9D",  -- 157
        66835 => X"87",  -- 135
        66836 => X"82",  -- 130
        66837 => X"9D",  -- 157
        66838 => X"9A",  -- 154
        66839 => X"95",  -- 149
        66840 => X"97",  -- 151
        66841 => X"B1",  -- 177
        66842 => X"A4",  -- 164
        66843 => X"9C",  -- 156
        66844 => X"98",  -- 152
        66845 => X"A8",  -- 168
        66846 => X"9B",  -- 155
        66847 => X"9D",  -- 157
        66848 => X"A1",  -- 161
        66849 => X"92",  -- 146
        66850 => X"8D",  -- 141
        66851 => X"98",  -- 152
        66852 => X"9A",  -- 154
        66853 => X"90",  -- 144
        66854 => X"89",  -- 137
        66855 => X"8E",  -- 142
        66856 => X"8A",  -- 138
        66857 => X"94",  -- 148
        66858 => X"97",  -- 151
        66859 => X"95",  -- 149
        66860 => X"A1",  -- 161
        66861 => X"B5",  -- 181
        66862 => X"B6",  -- 182
        66863 => X"AB",  -- 171
        66864 => X"A8",  -- 168
        66865 => X"A1",  -- 161
        66866 => X"8B",  -- 139
        66867 => X"96",  -- 150
        66868 => X"96",  -- 150
        66869 => X"A1",  -- 161
        66870 => X"9A",  -- 154
        66871 => X"A8",  -- 168
        66872 => X"A6",  -- 166
        66873 => X"B3",  -- 179
        66874 => X"B5",  -- 181
        66875 => X"A1",  -- 161
        66876 => X"9C",  -- 156
        66877 => X"9B",  -- 155
        66878 => X"97",  -- 151
        66879 => X"AC",  -- 172
        66880 => X"71",  -- 113
        66881 => X"77",  -- 119
        66882 => X"74",  -- 116
        66883 => X"6B",  -- 107
        66884 => X"6B",  -- 107
        66885 => X"6A",  -- 106
        66886 => X"5E",  -- 94
        66887 => X"57",  -- 87
        66888 => X"50",  -- 80
        66889 => X"52",  -- 82
        66890 => X"4F",  -- 79
        66891 => X"52",  -- 82
        66892 => X"54",  -- 84
        66893 => X"48",  -- 72
        66894 => X"38",  -- 56
        66895 => X"37",  -- 55
        66896 => X"4F",  -- 79
        66897 => X"67",  -- 103
        66898 => X"58",  -- 88
        66899 => X"4C",  -- 76
        66900 => X"55",  -- 85
        66901 => X"50",  -- 80
        66902 => X"47",  -- 71
        66903 => X"50",  -- 80
        66904 => X"49",  -- 73
        66905 => X"5B",  -- 91
        66906 => X"65",  -- 101
        66907 => X"73",  -- 115
        66908 => X"74",  -- 116
        66909 => X"52",  -- 82
        66910 => X"64",  -- 100
        66911 => X"67",  -- 103
        66912 => X"51",  -- 81
        66913 => X"55",  -- 85
        66914 => X"69",  -- 105
        66915 => X"4E",  -- 78
        66916 => X"81",  -- 129
        66917 => X"61",  -- 97
        66918 => X"5E",  -- 94
        66919 => X"7F",  -- 127
        66920 => X"69",  -- 105
        66921 => X"4D",  -- 77
        66922 => X"6B",  -- 107
        66923 => X"5C",  -- 92
        66924 => X"53",  -- 83
        66925 => X"8D",  -- 141
        66926 => X"7F",  -- 127
        66927 => X"4F",  -- 79
        66928 => X"59",  -- 89
        66929 => X"73",  -- 115
        66930 => X"79",  -- 121
        66931 => X"47",  -- 71
        66932 => X"52",  -- 82
        66933 => X"6A",  -- 106
        66934 => X"54",  -- 84
        66935 => X"59",  -- 89
        66936 => X"4C",  -- 76
        66937 => X"60",  -- 96
        66938 => X"4A",  -- 74
        66939 => X"45",  -- 69
        66940 => X"52",  -- 82
        66941 => X"4D",  -- 77
        66942 => X"4C",  -- 76
        66943 => X"4C",  -- 76
        66944 => X"46",  -- 70
        66945 => X"49",  -- 73
        66946 => X"50",  -- 80
        66947 => X"52",  -- 82
        66948 => X"4C",  -- 76
        66949 => X"45",  -- 69
        66950 => X"47",  -- 71
        66951 => X"4B",  -- 75
        66952 => X"4C",  -- 76
        66953 => X"36",  -- 54
        66954 => X"23",  -- 35
        66955 => X"34",  -- 52
        66956 => X"31",  -- 49
        66957 => X"3D",  -- 61
        66958 => X"5B",  -- 91
        66959 => X"4F",  -- 79
        66960 => X"42",  -- 66
        66961 => X"33",  -- 51
        66962 => X"4D",  -- 77
        66963 => X"5C",  -- 92
        66964 => X"67",  -- 103
        66965 => X"51",  -- 81
        66966 => X"4B",  -- 75
        66967 => X"82",  -- 130
        66968 => X"64",  -- 100
        66969 => X"58",  -- 88
        66970 => X"77",  -- 119
        66971 => X"5C",  -- 92
        66972 => X"24",  -- 36
        66973 => X"2B",  -- 43
        66974 => X"50",  -- 80
        66975 => X"4B",  -- 75
        66976 => X"37",  -- 55
        66977 => X"41",  -- 65
        66978 => X"6E",  -- 110
        66979 => X"8D",  -- 141
        66980 => X"72",  -- 114
        66981 => X"54",  -- 84
        66982 => X"2C",  -- 44
        66983 => X"4F",  -- 79
        66984 => X"8A",  -- 138
        66985 => X"69",  -- 105
        66986 => X"2D",  -- 45
        66987 => X"4B",  -- 75
        66988 => X"62",  -- 98
        66989 => X"5F",  -- 95
        66990 => X"50",  -- 80
        66991 => X"58",  -- 88
        66992 => X"73",  -- 115
        66993 => X"5D",  -- 93
        66994 => X"5C",  -- 92
        66995 => X"67",  -- 103
        66996 => X"61",  -- 97
        66997 => X"53",  -- 83
        66998 => X"4C",  -- 76
        66999 => X"47",  -- 71
        67000 => X"3C",  -- 60
        67001 => X"3A",  -- 58
        67002 => X"3D",  -- 61
        67003 => X"45",  -- 69
        67004 => X"45",  -- 69
        67005 => X"3B",  -- 59
        67006 => X"36",  -- 54
        67007 => X"36",  -- 54
        67008 => X"28",  -- 40
        67009 => X"24",  -- 36
        67010 => X"45",  -- 69
        67011 => X"55",  -- 85
        67012 => X"72",  -- 114
        67013 => X"68",  -- 104
        67014 => X"55",  -- 85
        67015 => X"56",  -- 86
        67016 => X"5D",  -- 93
        67017 => X"65",  -- 101
        67018 => X"5E",  -- 94
        67019 => X"5D",  -- 93
        67020 => X"80",  -- 128
        67021 => X"5F",  -- 95
        67022 => X"20",  -- 32
        67023 => X"12",  -- 18
        67024 => X"0A",  -- 10
        67025 => X"25",  -- 37
        67026 => X"35",  -- 53
        67027 => X"13",  -- 19
        67028 => X"3C",  -- 60
        67029 => X"00",  -- 0
        67030 => X"0C",  -- 12
        67031 => X"13",  -- 19
        67032 => X"3E",  -- 62
        67033 => X"4F",  -- 79
        67034 => X"4A",  -- 74
        67035 => X"1B",  -- 27
        67036 => X"0C",  -- 12
        67037 => X"27",  -- 39
        67038 => X"28",  -- 40
        67039 => X"1A",  -- 26
        67040 => X"5A",  -- 90
        67041 => X"2E",  -- 46
        67042 => X"29",  -- 41
        67043 => X"3D",  -- 61
        67044 => X"67",  -- 103
        67045 => X"2A",  -- 42
        67046 => X"36",  -- 54
        67047 => X"30",  -- 48
        67048 => X"2D",  -- 45
        67049 => X"2B",  -- 43
        67050 => X"29",  -- 41
        67051 => X"2D",  -- 45
        67052 => X"33",  -- 51
        67053 => X"37",  -- 55
        67054 => X"38",  -- 56
        67055 => X"38",  -- 56
        67056 => X"32",  -- 50
        67057 => X"3A",  -- 58
        67058 => X"3B",  -- 59
        67059 => X"39",  -- 57
        67060 => X"3B",  -- 59
        67061 => X"39",  -- 57
        67062 => X"3B",  -- 59
        67063 => X"44",  -- 68
        67064 => X"42",  -- 66
        67065 => X"3F",  -- 63
        67066 => X"42",  -- 66
        67067 => X"48",  -- 72
        67068 => X"4A",  -- 74
        67069 => X"49",  -- 73
        67070 => X"4B",  -- 75
        67071 => X"50",  -- 80
        67072 => X"4B",  -- 75
        67073 => X"4D",  -- 77
        67074 => X"50",  -- 80
        67075 => X"57",  -- 87
        67076 => X"5B",  -- 91
        67077 => X"5E",  -- 94
        67078 => X"67",  -- 103
        67079 => X"70",  -- 112
        67080 => X"70",  -- 112
        67081 => X"71",  -- 113
        67082 => X"66",  -- 102
        67083 => X"62",  -- 98
        67084 => X"65",  -- 101
        67085 => X"56",  -- 86
        67086 => X"41",  -- 65
        67087 => X"3F",  -- 63
        67088 => X"53",  -- 83
        67089 => X"56",  -- 86
        67090 => X"4F",  -- 79
        67091 => X"42",  -- 66
        67092 => X"37",  -- 55
        67093 => X"34",  -- 52
        67094 => X"2F",  -- 47
        67095 => X"26",  -- 38
        67096 => X"27",  -- 39
        67097 => X"22",  -- 34
        67098 => X"15",  -- 21
        67099 => X"08",  -- 8
        67100 => X"07",  -- 7
        67101 => X"12",  -- 18
        67102 => X"1D",  -- 29
        67103 => X"24",  -- 36
        67104 => X"45",  -- 69
        67105 => X"5C",  -- 92
        67106 => X"67",  -- 103
        67107 => X"6B",  -- 107
        67108 => X"7B",  -- 123
        67109 => X"75",  -- 117
        67110 => X"62",  -- 98
        67111 => X"6A",  -- 106
        67112 => X"7B",  -- 123
        67113 => X"95",  -- 149
        67114 => X"A9",  -- 169
        67115 => X"A3",  -- 163
        67116 => X"8F",  -- 143
        67117 => X"87",  -- 135
        67118 => X"8E",  -- 142
        67119 => X"97",  -- 151
        67120 => X"93",  -- 147
        67121 => X"92",  -- 146
        67122 => X"8A",  -- 138
        67123 => X"8B",  -- 139
        67124 => X"8C",  -- 140
        67125 => X"8F",  -- 143
        67126 => X"9D",  -- 157
        67127 => X"9E",  -- 158
        67128 => X"8D",  -- 141
        67129 => X"8A",  -- 138
        67130 => X"96",  -- 150
        67131 => X"9F",  -- 159
        67132 => X"93",  -- 147
        67133 => X"82",  -- 130
        67134 => X"80",  -- 128
        67135 => X"85",  -- 133
        67136 => X"88",  -- 136
        67137 => X"85",  -- 133
        67138 => X"88",  -- 136
        67139 => X"8C",  -- 140
        67140 => X"8D",  -- 141
        67141 => X"96",  -- 150
        67142 => X"9F",  -- 159
        67143 => X"9F",  -- 159
        67144 => X"96",  -- 150
        67145 => X"9B",  -- 155
        67146 => X"9F",  -- 159
        67147 => X"94",  -- 148
        67148 => X"93",  -- 147
        67149 => X"95",  -- 149
        67150 => X"A3",  -- 163
        67151 => X"A7",  -- 167
        67152 => X"96",  -- 150
        67153 => X"9A",  -- 154
        67154 => X"A2",  -- 162
        67155 => X"A0",  -- 160
        67156 => X"90",  -- 144
        67157 => X"93",  -- 147
        67158 => X"A3",  -- 163
        67159 => X"9D",  -- 157
        67160 => X"79",  -- 121
        67161 => X"8A",  -- 138
        67162 => X"8A",  -- 138
        67163 => X"93",  -- 147
        67164 => X"A0",  -- 160
        67165 => X"A5",  -- 165
        67166 => X"96",  -- 150
        67167 => X"93",  -- 147
        67168 => X"8A",  -- 138
        67169 => X"9F",  -- 159
        67170 => X"A0",  -- 160
        67171 => X"8D",  -- 141
        67172 => X"8F",  -- 143
        67173 => X"A5",  -- 165
        67174 => X"A5",  -- 165
        67175 => X"8F",  -- 143
        67176 => X"9A",  -- 154
        67177 => X"9B",  -- 155
        67178 => X"98",  -- 152
        67179 => X"95",  -- 149
        67180 => X"97",  -- 151
        67181 => X"A0",  -- 160
        67182 => X"AA",  -- 170
        67183 => X"B0",  -- 176
        67184 => X"93",  -- 147
        67185 => X"98",  -- 152
        67186 => X"90",  -- 144
        67187 => X"A0",  -- 160
        67188 => X"A5",  -- 165
        67189 => X"AD",  -- 173
        67190 => X"A1",  -- 161
        67191 => X"A7",  -- 167
        67192 => X"BD",  -- 189
        67193 => X"B3",  -- 179
        67194 => X"A9",  -- 169
        67195 => X"97",  -- 151
        67196 => X"9A",  -- 154
        67197 => X"A5",  -- 165
        67198 => X"A2",  -- 162
        67199 => X"AB",  -- 171
        67200 => X"76",  -- 118
        67201 => X"79",  -- 121
        67202 => X"79",  -- 121
        67203 => X"72",  -- 114
        67204 => X"68",  -- 104
        67205 => X"6A",  -- 106
        67206 => X"6A",  -- 106
        67207 => X"62",  -- 98
        67208 => X"52",  -- 82
        67209 => X"5B",  -- 91
        67210 => X"66",  -- 102
        67211 => X"6F",  -- 111
        67212 => X"6B",  -- 107
        67213 => X"52",  -- 82
        67214 => X"40",  -- 64
        67215 => X"42",  -- 66
        67216 => X"5E",  -- 94
        67217 => X"7F",  -- 127
        67218 => X"5D",  -- 93
        67219 => X"5F",  -- 95
        67220 => X"7B",  -- 123
        67221 => X"61",  -- 97
        67222 => X"51",  -- 81
        67223 => X"56",  -- 86
        67224 => X"62",  -- 98
        67225 => X"66",  -- 102
        67226 => X"6A",  -- 106
        67227 => X"71",  -- 113
        67228 => X"6B",  -- 107
        67229 => X"56",  -- 86
        67230 => X"6D",  -- 109
        67231 => X"5C",  -- 92
        67232 => X"56",  -- 86
        67233 => X"6E",  -- 110
        67234 => X"66",  -- 102
        67235 => X"6A",  -- 106
        67236 => X"88",  -- 136
        67237 => X"4A",  -- 74
        67238 => X"5E",  -- 94
        67239 => X"83",  -- 131
        67240 => X"5D",  -- 93
        67241 => X"51",  -- 81
        67242 => X"77",  -- 119
        67243 => X"51",  -- 81
        67244 => X"66",  -- 102
        67245 => X"9A",  -- 154
        67246 => X"61",  -- 97
        67247 => X"4F",  -- 79
        67248 => X"6A",  -- 106
        67249 => X"86",  -- 134
        67250 => X"69",  -- 105
        67251 => X"3E",  -- 62
        67252 => X"65",  -- 101
        67253 => X"5C",  -- 92
        67254 => X"54",  -- 84
        67255 => X"57",  -- 87
        67256 => X"52",  -- 82
        67257 => X"5D",  -- 93
        67258 => X"47",  -- 71
        67259 => X"41",  -- 65
        67260 => X"50",  -- 80
        67261 => X"4F",  -- 79
        67262 => X"4C",  -- 76
        67263 => X"4B",  -- 75
        67264 => X"4C",  -- 76
        67265 => X"49",  -- 73
        67266 => X"48",  -- 72
        67267 => X"4A",  -- 74
        67268 => X"49",  -- 73
        67269 => X"47",  -- 71
        67270 => X"49",  -- 73
        67271 => X"4C",  -- 76
        67272 => X"3F",  -- 63
        67273 => X"2E",  -- 46
        67274 => X"20",  -- 32
        67275 => X"2F",  -- 47
        67276 => X"2A",  -- 42
        67277 => X"55",  -- 85
        67278 => X"5A",  -- 90
        67279 => X"3F",  -- 63
        67280 => X"49",  -- 73
        67281 => X"39",  -- 57
        67282 => X"45",  -- 69
        67283 => X"53",  -- 83
        67284 => X"66",  -- 102
        67285 => X"3E",  -- 62
        67286 => X"47",  -- 71
        67287 => X"6F",  -- 111
        67288 => X"3C",  -- 60
        67289 => X"3E",  -- 62
        67290 => X"7C",  -- 124
        67291 => X"5E",  -- 94
        67292 => X"21",  -- 33
        67293 => X"1E",  -- 30
        67294 => X"48",  -- 72
        67295 => X"35",  -- 53
        67296 => X"35",  -- 53
        67297 => X"3F",  -- 63
        67298 => X"55",  -- 85
        67299 => X"92",  -- 146
        67300 => X"60",  -- 96
        67301 => X"41",  -- 65
        67302 => X"2C",  -- 44
        67303 => X"30",  -- 48
        67304 => X"80",  -- 128
        67305 => X"54",  -- 84
        67306 => X"35",  -- 53
        67307 => X"2F",  -- 47
        67308 => X"48",  -- 72
        67309 => X"50",  -- 80
        67310 => X"63",  -- 99
        67311 => X"50",  -- 80
        67312 => X"66",  -- 102
        67313 => X"5D",  -- 93
        67314 => X"4E",  -- 78
        67315 => X"58",  -- 88
        67316 => X"6C",  -- 108
        67317 => X"59",  -- 89
        67318 => X"41",  -- 65
        67319 => X"4D",  -- 77
        67320 => X"3D",  -- 61
        67321 => X"3B",  -- 59
        67322 => X"3B",  -- 59
        67323 => X"3C",  -- 60
        67324 => X"3E",  -- 62
        67325 => X"3F",  -- 63
        67326 => X"3D",  -- 61
        67327 => X"3A",  -- 58
        67328 => X"39",  -- 57
        67329 => X"19",  -- 25
        67330 => X"3A",  -- 58
        67331 => X"42",  -- 66
        67332 => X"5F",  -- 95
        67333 => X"6C",  -- 108
        67334 => X"57",  -- 87
        67335 => X"5B",  -- 91
        67336 => X"5B",  -- 91
        67337 => X"66",  -- 102
        67338 => X"52",  -- 82
        67339 => X"4F",  -- 79
        67340 => X"7B",  -- 123
        67341 => X"67",  -- 103
        67342 => X"10",  -- 16
        67343 => X"0C",  -- 12
        67344 => X"02",  -- 2
        67345 => X"0A",  -- 10
        67346 => X"49",  -- 73
        67347 => X"07",  -- 7
        67348 => X"46",  -- 70
        67349 => X"1B",  -- 27
        67350 => X"08",  -- 8
        67351 => X"10",  -- 16
        67352 => X"12",  -- 18
        67353 => X"0E",  -- 14
        67354 => X"35",  -- 53
        67355 => X"57",  -- 87
        67356 => X"4C",  -- 76
        67357 => X"22",  -- 34
        67358 => X"16",  -- 22
        67359 => X"39",  -- 57
        67360 => X"4E",  -- 78
        67361 => X"57",  -- 87
        67362 => X"1F",  -- 31
        67363 => X"1A",  -- 26
        67364 => X"50",  -- 80
        67365 => X"4F",  -- 79
        67366 => X"22",  -- 34
        67367 => X"2B",  -- 43
        67368 => X"2C",  -- 44
        67369 => X"2C",  -- 44
        67370 => X"2A",  -- 42
        67371 => X"2D",  -- 45
        67372 => X"33",  -- 51
        67373 => X"39",  -- 57
        67374 => X"3B",  -- 59
        67375 => X"38",  -- 56
        67376 => X"2D",  -- 45
        67377 => X"39",  -- 57
        67378 => X"3D",  -- 61
        67379 => X"40",  -- 64
        67380 => X"46",  -- 70
        67381 => X"46",  -- 70
        67382 => X"48",  -- 72
        67383 => X"4F",  -- 79
        67384 => X"4E",  -- 78
        67385 => X"4B",  -- 75
        67386 => X"4E",  -- 78
        67387 => X"55",  -- 85
        67388 => X"4F",  -- 79
        67389 => X"45",  -- 69
        67390 => X"4B",  -- 75
        67391 => X"5C",  -- 92
        67392 => X"56",  -- 86
        67393 => X"57",  -- 87
        67394 => X"59",  -- 89
        67395 => X"5D",  -- 93
        67396 => X"5E",  -- 94
        67397 => X"5F",  -- 95
        67398 => X"68",  -- 104
        67399 => X"70",  -- 112
        67400 => X"74",  -- 116
        67401 => X"72",  -- 114
        67402 => X"68",  -- 104
        67403 => X"62",  -- 98
        67404 => X"62",  -- 98
        67405 => X"54",  -- 84
        67406 => X"45",  -- 69
        67407 => X"44",  -- 68
        67408 => X"4D",  -- 77
        67409 => X"48",  -- 72
        67410 => X"3C",  -- 60
        67411 => X"2F",  -- 47
        67412 => X"2C",  -- 44
        67413 => X"2D",  -- 45
        67414 => X"2A",  -- 42
        67415 => X"20",  -- 32
        67416 => X"15",  -- 21
        67417 => X"15",  -- 21
        67418 => X"10",  -- 16
        67419 => X"07",  -- 7
        67420 => X"02",  -- 2
        67421 => X"05",  -- 5
        67422 => X"0C",  -- 12
        67423 => X"10",  -- 16
        67424 => X"31",  -- 49
        67425 => X"49",  -- 73
        67426 => X"51",  -- 81
        67427 => X"59",  -- 89
        67428 => X"6F",  -- 111
        67429 => X"73",  -- 115
        67430 => X"68",  -- 104
        67431 => X"63",  -- 99
        67432 => X"79",  -- 121
        67433 => X"89",  -- 137
        67434 => X"94",  -- 148
        67435 => X"93",  -- 147
        67436 => X"92",  -- 146
        67437 => X"98",  -- 152
        67438 => X"9C",  -- 156
        67439 => X"98",  -- 152
        67440 => X"96",  -- 150
        67441 => X"85",  -- 133
        67442 => X"8C",  -- 140
        67443 => X"8E",  -- 142
        67444 => X"8E",  -- 142
        67445 => X"9E",  -- 158
        67446 => X"A3",  -- 163
        67447 => X"A0",  -- 160
        67448 => X"95",  -- 149
        67449 => X"93",  -- 147
        67450 => X"93",  -- 147
        67451 => X"92",  -- 146
        67452 => X"8E",  -- 142
        67453 => X"89",  -- 137
        67454 => X"88",  -- 136
        67455 => X"89",  -- 137
        67456 => X"95",  -- 149
        67457 => X"97",  -- 151
        67458 => X"92",  -- 146
        67459 => X"8F",  -- 143
        67460 => X"93",  -- 147
        67461 => X"95",  -- 149
        67462 => X"97",  -- 151
        67463 => X"9D",  -- 157
        67464 => X"98",  -- 152
        67465 => X"A1",  -- 161
        67466 => X"97",  -- 151
        67467 => X"86",  -- 134
        67468 => X"79",  -- 121
        67469 => X"88",  -- 136
        67470 => X"8F",  -- 143
        67471 => X"90",  -- 144
        67472 => X"91",  -- 145
        67473 => X"94",  -- 148
        67474 => X"97",  -- 151
        67475 => X"A6",  -- 166
        67476 => X"8C",  -- 140
        67477 => X"77",  -- 119
        67478 => X"87",  -- 135
        67479 => X"70",  -- 112
        67480 => X"8F",  -- 143
        67481 => X"94",  -- 148
        67482 => X"99",  -- 153
        67483 => X"9B",  -- 155
        67484 => X"A7",  -- 167
        67485 => X"9E",  -- 158
        67486 => X"9C",  -- 156
        67487 => X"9F",  -- 159
        67488 => X"98",  -- 152
        67489 => X"A0",  -- 160
        67490 => X"A2",  -- 162
        67491 => X"9C",  -- 156
        67492 => X"9A",  -- 154
        67493 => X"A0",  -- 160
        67494 => X"A1",  -- 161
        67495 => X"9C",  -- 156
        67496 => X"AA",  -- 170
        67497 => X"AD",  -- 173
        67498 => X"B5",  -- 181
        67499 => X"BA",  -- 186
        67500 => X"B2",  -- 178
        67501 => X"A5",  -- 165
        67502 => X"A5",  -- 165
        67503 => X"AE",  -- 174
        67504 => X"A6",  -- 166
        67505 => X"AD",  -- 173
        67506 => X"A6",  -- 166
        67507 => X"A9",  -- 169
        67508 => X"A9",  -- 169
        67509 => X"AA",  -- 170
        67510 => X"99",  -- 153
        67511 => X"95",  -- 149
        67512 => X"82",  -- 130
        67513 => X"81",  -- 129
        67514 => X"8F",  -- 143
        67515 => X"8B",  -- 139
        67516 => X"86",  -- 134
        67517 => X"8D",  -- 141
        67518 => X"89",  -- 137
        67519 => X"8A",  -- 138
        67520 => X"7A",  -- 122
        67521 => X"77",  -- 119
        67522 => X"7D",  -- 125
        67523 => X"78",  -- 120
        67524 => X"6D",  -- 109
        67525 => X"75",  -- 117
        67526 => X"7D",  -- 125
        67527 => X"73",  -- 115
        67528 => X"63",  -- 99
        67529 => X"69",  -- 105
        67530 => X"70",  -- 112
        67531 => X"79",  -- 121
        67532 => X"75",  -- 117
        67533 => X"61",  -- 97
        67534 => X"58",  -- 88
        67535 => X"63",  -- 99
        67536 => X"7A",  -- 122
        67537 => X"70",  -- 112
        67538 => X"65",  -- 101
        67539 => X"72",  -- 114
        67540 => X"6F",  -- 111
        67541 => X"63",  -- 99
        67542 => X"63",  -- 99
        67543 => X"52",  -- 82
        67544 => X"6C",  -- 108
        67545 => X"61",  -- 97
        67546 => X"63",  -- 99
        67547 => X"6A",  -- 106
        67548 => X"69",  -- 105
        67549 => X"66",  -- 102
        67550 => X"80",  -- 128
        67551 => X"5C",  -- 92
        67552 => X"5D",  -- 93
        67553 => X"77",  -- 119
        67554 => X"61",  -- 97
        67555 => X"8D",  -- 141
        67556 => X"63",  -- 99
        67557 => X"5A",  -- 90
        67558 => X"54",  -- 84
        67559 => X"8C",  -- 140
        67560 => X"59",  -- 89
        67561 => X"5D",  -- 93
        67562 => X"81",  -- 129
        67563 => X"50",  -- 80
        67564 => X"7E",  -- 126
        67565 => X"88",  -- 136
        67566 => X"4E",  -- 78
        67567 => X"5A",  -- 90
        67568 => X"84",  -- 132
        67569 => X"8C",  -- 140
        67570 => X"58",  -- 88
        67571 => X"4D",  -- 77
        67572 => X"6A",  -- 106
        67573 => X"50",  -- 80
        67574 => X"54",  -- 84
        67575 => X"51",  -- 81
        67576 => X"52",  -- 82
        67577 => X"59",  -- 89
        67578 => X"4B",  -- 75
        67579 => X"46",  -- 70
        67580 => X"4E",  -- 78
        67581 => X"4F",  -- 79
        67582 => X"4B",  -- 75
        67583 => X"4B",  -- 75
        67584 => X"54",  -- 84
        67585 => X"45",  -- 69
        67586 => X"3B",  -- 59
        67587 => X"42",  -- 66
        67588 => X"4D",  -- 77
        67589 => X"50",  -- 80
        67590 => X"49",  -- 73
        67591 => X"40",  -- 64
        67592 => X"35",  -- 53
        67593 => X"37",  -- 55
        67594 => X"34",  -- 52
        67595 => X"38",  -- 56
        67596 => X"49",  -- 73
        67597 => X"6A",  -- 106
        67598 => X"50",  -- 80
        67599 => X"34",  -- 52
        67600 => X"41",  -- 65
        67601 => X"38",  -- 56
        67602 => X"3E",  -- 62
        67603 => X"50",  -- 80
        67604 => X"6A",  -- 106
        67605 => X"32",  -- 50
        67606 => X"3F",  -- 63
        67607 => X"52",  -- 82
        67608 => X"2E",  -- 46
        67609 => X"2F",  -- 47
        67610 => X"65",  -- 101
        67611 => X"4A",  -- 74
        67612 => X"31",  -- 49
        67613 => X"24",  -- 36
        67614 => X"3A",  -- 58
        67615 => X"25",  -- 37
        67616 => X"39",  -- 57
        67617 => X"39",  -- 57
        67618 => X"4F",  -- 79
        67619 => X"7D",  -- 125
        67620 => X"4B",  -- 75
        67621 => X"3D",  -- 61
        67622 => X"38",  -- 56
        67623 => X"26",  -- 38
        67624 => X"6F",  -- 111
        67625 => X"44",  -- 68
        67626 => X"42",  -- 66
        67627 => X"36",  -- 54
        67628 => X"3E",  -- 62
        67629 => X"4A",  -- 74
        67630 => X"6A",  -- 106
        67631 => X"4C",  -- 76
        67632 => X"5E",  -- 94
        67633 => X"59",  -- 89
        67634 => X"48",  -- 72
        67635 => X"4E",  -- 78
        67636 => X"64",  -- 100
        67637 => X"59",  -- 89
        67638 => X"41",  -- 65
        67639 => X"42",  -- 66
        67640 => X"3D",  -- 61
        67641 => X"3B",  -- 59
        67642 => X"36",  -- 54
        67643 => X"31",  -- 49
        67644 => X"35",  -- 53
        67645 => X"3E",  -- 62
        67646 => X"3F",  -- 63
        67647 => X"3A",  -- 58
        67648 => X"4B",  -- 75
        67649 => X"23",  -- 35
        67650 => X"2F",  -- 47
        67651 => X"38",  -- 56
        67652 => X"4A",  -- 74
        67653 => X"61",  -- 97
        67654 => X"5C",  -- 92
        67655 => X"5F",  -- 95
        67656 => X"4C",  -- 76
        67657 => X"57",  -- 87
        67658 => X"48",  -- 72
        67659 => X"41",  -- 65
        67660 => X"5E",  -- 94
        67661 => X"66",  -- 102
        67662 => X"14",  -- 20
        67663 => X"02",  -- 2
        67664 => X"09",  -- 9
        67665 => X"04",  -- 4
        67666 => X"34",  -- 52
        67667 => X"17",  -- 23
        67668 => X"28",  -- 40
        67669 => X"3E",  -- 62
        67670 => X"14",  -- 20
        67671 => X"14",  -- 20
        67672 => X"1B",  -- 27
        67673 => X"0D",  -- 13
        67674 => X"0B",  -- 11
        67675 => X"10",  -- 16
        67676 => X"34",  -- 52
        67677 => X"55",  -- 85
        67678 => X"43",  -- 67
        67679 => X"29",  -- 41
        67680 => X"2B",  -- 43
        67681 => X"55",  -- 85
        67682 => X"1D",  -- 29
        67683 => X"1C",  -- 28
        67684 => X"32",  -- 50
        67685 => X"6F",  -- 111
        67686 => X"33",  -- 51
        67687 => X"38",  -- 56
        67688 => X"27",  -- 39
        67689 => X"31",  -- 49
        67690 => X"39",  -- 57
        67691 => X"39",  -- 57
        67692 => X"37",  -- 55
        67693 => X"38",  -- 56
        67694 => X"3A",  -- 58
        67695 => X"3C",  -- 60
        67696 => X"3F",  -- 63
        67697 => X"40",  -- 64
        67698 => X"3E",  -- 62
        67699 => X"42",  -- 66
        67700 => X"51",  -- 81
        67701 => X"57",  -- 87
        67702 => X"53",  -- 83
        67703 => X"55",  -- 85
        67704 => X"55",  -- 85
        67705 => X"56",  -- 86
        67706 => X"59",  -- 89
        67707 => X"59",  -- 89
        67708 => X"52",  -- 82
        67709 => X"4C",  -- 76
        67710 => X"54",  -- 84
        67711 => X"61",  -- 97
        67712 => X"59",  -- 89
        67713 => X"5B",  -- 91
        67714 => X"5D",  -- 93
        67715 => X"61",  -- 97
        67716 => X"5F",  -- 95
        67717 => X"5E",  -- 94
        67718 => X"64",  -- 100
        67719 => X"6B",  -- 107
        67720 => X"75",  -- 117
        67721 => X"70",  -- 112
        67722 => X"69",  -- 105
        67723 => X"65",  -- 101
        67724 => X"5F",  -- 95
        67725 => X"52",  -- 82
        67726 => X"4A",  -- 74
        67727 => X"4A",  -- 74
        67728 => X"44",  -- 68
        67729 => X"3D",  -- 61
        67730 => X"2F",  -- 47
        67731 => X"22",  -- 34
        67732 => X"22",  -- 34
        67733 => X"25",  -- 37
        67734 => X"25",  -- 37
        67735 => X"1E",  -- 30
        67736 => X"11",  -- 17
        67737 => X"12",  -- 18
        67738 => X"10",  -- 16
        67739 => X"0C",  -- 12
        67740 => X"09",  -- 9
        67741 => X"09",  -- 9
        67742 => X"0B",  -- 11
        67743 => X"0C",  -- 12
        67744 => X"12",  -- 18
        67745 => X"22",  -- 34
        67746 => X"24",  -- 36
        67747 => X"35",  -- 53
        67748 => X"54",  -- 84
        67749 => X"62",  -- 98
        67750 => X"68",  -- 104
        67751 => X"6A",  -- 106
        67752 => X"81",  -- 129
        67753 => X"8B",  -- 139
        67754 => X"8D",  -- 141
        67755 => X"83",  -- 131
        67756 => X"80",  -- 128
        67757 => X"8C",  -- 140
        67758 => X"92",  -- 146
        67759 => X"90",  -- 144
        67760 => X"99",  -- 153
        67761 => X"81",  -- 129
        67762 => X"94",  -- 148
        67763 => X"94",  -- 148
        67764 => X"8C",  -- 140
        67765 => X"9B",  -- 155
        67766 => X"95",  -- 149
        67767 => X"8C",  -- 140
        67768 => X"97",  -- 151
        67769 => X"97",  -- 151
        67770 => X"8A",  -- 138
        67771 => X"81",  -- 129
        67772 => X"91",  -- 145
        67773 => X"A2",  -- 162
        67774 => X"9C",  -- 156
        67775 => X"8E",  -- 142
        67776 => X"87",  -- 135
        67777 => X"91",  -- 145
        67778 => X"8D",  -- 141
        67779 => X"8E",  -- 142
        67780 => X"9B",  -- 155
        67781 => X"9D",  -- 157
        67782 => X"9A",  -- 154
        67783 => X"A4",  -- 164
        67784 => X"A8",  -- 168
        67785 => X"A5",  -- 165
        67786 => X"8E",  -- 142
        67787 => X"8B",  -- 139
        67788 => X"86",  -- 134
        67789 => X"9C",  -- 156
        67790 => X"98",  -- 152
        67791 => X"95",  -- 149
        67792 => X"9A",  -- 154
        67793 => X"8A",  -- 138
        67794 => X"86",  -- 134
        67795 => X"92",  -- 146
        67796 => X"88",  -- 136
        67797 => X"8B",  -- 139
        67798 => X"9D",  -- 157
        67799 => X"87",  -- 135
        67800 => X"91",  -- 145
        67801 => X"8D",  -- 141
        67802 => X"8B",  -- 139
        67803 => X"74",  -- 116
        67804 => X"78",  -- 120
        67805 => X"7C",  -- 124
        67806 => X"A1",  -- 161
        67807 => X"BA",  -- 186
        67808 => X"B1",  -- 177
        67809 => X"A5",  -- 165
        67810 => X"A7",  -- 167
        67811 => X"B7",  -- 183
        67812 => X"B5",  -- 181
        67813 => X"A3",  -- 163
        67814 => X"A2",  -- 162
        67815 => X"B1",  -- 177
        67816 => X"BB",  -- 187
        67817 => X"B5",  -- 181
        67818 => X"B2",  -- 178
        67819 => X"B1",  -- 177
        67820 => X"AC",  -- 172
        67821 => X"A8",  -- 168
        67822 => X"AD",  -- 173
        67823 => X"B8",  -- 184
        67824 => X"AC",  -- 172
        67825 => X"AE",  -- 174
        67826 => X"9D",  -- 157
        67827 => X"8E",  -- 142
        67828 => X"8B",  -- 139
        67829 => X"8B",  -- 139
        67830 => X"83",  -- 131
        67831 => X"80",  -- 128
        67832 => X"8A",  -- 138
        67833 => X"82",  -- 130
        67834 => X"90",  -- 144
        67835 => X"8B",  -- 139
        67836 => X"83",  -- 131
        67837 => X"93",  -- 147
        67838 => X"9D",  -- 157
        67839 => X"A0",  -- 160
        67840 => X"7A",  -- 122
        67841 => X"77",  -- 119
        67842 => X"7A",  -- 122
        67843 => X"76",  -- 118
        67844 => X"6D",  -- 109
        67845 => X"77",  -- 119
        67846 => X"81",  -- 129
        67847 => X"76",  -- 118
        67848 => X"78",  -- 120
        67849 => X"75",  -- 117
        67850 => X"6F",  -- 111
        67851 => X"71",  -- 113
        67852 => X"73",  -- 115
        67853 => X"6B",  -- 107
        67854 => X"6C",  -- 108
        67855 => X"7C",  -- 124
        67856 => X"86",  -- 134
        67857 => X"60",  -- 96
        67858 => X"6C",  -- 108
        67859 => X"71",  -- 113
        67860 => X"5E",  -- 94
        67861 => X"69",  -- 105
        67862 => X"73",  -- 115
        67863 => X"6C",  -- 108
        67864 => X"73",  -- 115
        67865 => X"6A",  -- 106
        67866 => X"6F",  -- 111
        67867 => X"74",  -- 116
        67868 => X"6D",  -- 109
        67869 => X"69",  -- 105
        67870 => X"84",  -- 132
        67871 => X"57",  -- 87
        67872 => X"60",  -- 96
        67873 => X"5F",  -- 95
        67874 => X"75",  -- 117
        67875 => X"8A",  -- 138
        67876 => X"4D",  -- 77
        67877 => X"6B",  -- 107
        67878 => X"57",  -- 87
        67879 => X"88",  -- 136
        67880 => X"5C",  -- 92
        67881 => X"62",  -- 98
        67882 => X"75",  -- 117
        67883 => X"5C",  -- 92
        67884 => X"98",  -- 152
        67885 => X"71",  -- 113
        67886 => X"4E",  -- 78
        67887 => X"63",  -- 99
        67888 => X"92",  -- 146
        67889 => X"79",  -- 121
        67890 => X"4B",  -- 75
        67891 => X"64",  -- 100
        67892 => X"5F",  -- 95
        67893 => X"4D",  -- 77
        67894 => X"56",  -- 86
        67895 => X"4E",  -- 78
        67896 => X"4A",  -- 74
        67897 => X"4F",  -- 79
        67898 => X"52",  -- 82
        67899 => X"4F",  -- 79
        67900 => X"52",  -- 82
        67901 => X"53",  -- 83
        67902 => X"4E",  -- 78
        67903 => X"51",  -- 81
        67904 => X"53",  -- 83
        67905 => X"45",  -- 69
        67906 => X"3D",  -- 61
        67907 => X"45",  -- 69
        67908 => X"50",  -- 80
        67909 => X"51",  -- 81
        67910 => X"46",  -- 70
        67911 => X"3A",  -- 58
        67912 => X"3B",  -- 59
        67913 => X"3B",  -- 59
        67914 => X"3E",  -- 62
        67915 => X"47",  -- 71
        67916 => X"71",  -- 113
        67917 => X"5A",  -- 90
        67918 => X"33",  -- 51
        67919 => X"39",  -- 57
        67920 => X"32",  -- 50
        67921 => X"31",  -- 49
        67922 => X"33",  -- 51
        67923 => X"44",  -- 68
        67924 => X"60",  -- 96
        67925 => X"27",  -- 39
        67926 => X"34",  -- 52
        67927 => X"39",  -- 57
        67928 => X"2F",  -- 47
        67929 => X"2E",  -- 46
        67930 => X"48",  -- 72
        67931 => X"32",  -- 50
        67932 => X"40",  -- 64
        67933 => X"2B",  -- 43
        67934 => X"29",  -- 41
        67935 => X"25",  -- 37
        67936 => X"36",  -- 54
        67937 => X"2E",  -- 46
        67938 => X"56",  -- 86
        67939 => X"59",  -- 89
        67940 => X"39",  -- 57
        67941 => X"41",  -- 65
        67942 => X"3A",  -- 58
        67943 => X"20",  -- 32
        67944 => X"5D",  -- 93
        67945 => X"35",  -- 53
        67946 => X"3C",  -- 60
        67947 => X"39",  -- 57
        67948 => X"2A",  -- 42
        67949 => X"3B",  -- 59
        67950 => X"5E",  -- 94
        67951 => X"52",  -- 82
        67952 => X"5D",  -- 93
        67953 => X"54",  -- 84
        67954 => X"4B",  -- 75
        67955 => X"49",  -- 73
        67956 => X"4E",  -- 78
        67957 => X"54",  -- 84
        67958 => X"48",  -- 72
        67959 => X"2F",  -- 47
        67960 => X"34",  -- 52
        67961 => X"32",  -- 50
        67962 => X"2A",  -- 42
        67963 => X"21",  -- 33
        67964 => X"24",  -- 36
        67965 => X"30",  -- 48
        67966 => X"34",  -- 52
        67967 => X"2D",  -- 45
        67968 => X"3F",  -- 63
        67969 => X"29",  -- 41
        67970 => X"28",  -- 40
        67971 => X"3E",  -- 62
        67972 => X"44",  -- 68
        67973 => X"4D",  -- 77
        67974 => X"53",  -- 83
        67975 => X"4E",  -- 78
        67976 => X"48",  -- 72
        67977 => X"46",  -- 70
        67978 => X"42",  -- 66
        67979 => X"3E",  -- 62
        67980 => X"47",  -- 71
        67981 => X"6D",  -- 109
        67982 => X"3A",  -- 58
        67983 => X"01",  -- 1
        67984 => X"0F",  -- 15
        67985 => X"0D",  -- 13
        67986 => X"23",  -- 35
        67987 => X"3D",  -- 61
        67988 => X"12",  -- 18
        67989 => X"49",  -- 73
        67990 => X"30",  -- 48
        67991 => X"26",  -- 38
        67992 => X"30",  -- 48
        67993 => X"21",  -- 33
        67994 => X"23",  -- 35
        67995 => X"20",  -- 32
        67996 => X"1C",  -- 28
        67997 => X"1E",  -- 30
        67998 => X"26",  -- 38
        67999 => X"40",  -- 64
        68000 => X"4C",  -- 76
        68001 => X"5C",  -- 92
        68002 => X"6A",  -- 106
        68003 => X"3C",  -- 60
        68004 => X"41",  -- 65
        68005 => X"56",  -- 86
        68006 => X"53",  -- 83
        68007 => X"28",  -- 40
        68008 => X"36",  -- 54
        68009 => X"41",  -- 65
        68010 => X"49",  -- 73
        68011 => X"49",  -- 73
        68012 => X"45",  -- 69
        68013 => X"46",  -- 70
        68014 => X"48",  -- 72
        68015 => X"49",  -- 73
        68016 => X"4F",  -- 79
        68017 => X"51",  -- 81
        68018 => X"4E",  -- 78
        68019 => X"4F",  -- 79
        68020 => X"5A",  -- 90
        68021 => X"5B",  -- 91
        68022 => X"55",  -- 85
        68023 => X"55",  -- 85
        68024 => X"54",  -- 84
        68025 => X"5B",  -- 91
        68026 => X"5D",  -- 93
        68027 => X"58",  -- 88
        68028 => X"59",  -- 89
        68029 => X"5F",  -- 95
        68030 => X"65",  -- 101
        68031 => X"65",  -- 101
        68032 => X"5A",  -- 90
        68033 => X"5C",  -- 92
        68034 => X"60",  -- 96
        68035 => X"66",  -- 102
        68036 => X"66",  -- 102
        68037 => X"63",  -- 99
        68038 => X"63",  -- 99
        68039 => X"66",  -- 102
        68040 => X"6E",  -- 110
        68041 => X"68",  -- 104
        68042 => X"68",  -- 104
        68043 => X"65",  -- 101
        68044 => X"5C",  -- 92
        68045 => X"52",  -- 82
        68046 => X"4D",  -- 77
        68047 => X"4C",  -- 76
        68048 => X"45",  -- 69
        68049 => X"3D",  -- 61
        68050 => X"2F",  -- 47
        68051 => X"23",  -- 35
        68052 => X"1F",  -- 31
        68053 => X"20",  -- 32
        68054 => X"1E",  -- 30
        68055 => X"1C",  -- 28
        68056 => X"16",  -- 22
        68057 => X"12",  -- 18
        68058 => X"10",  -- 16
        68059 => X"11",  -- 17
        68060 => X"13",  -- 19
        68061 => X"14",  -- 20
        68062 => X"15",  -- 21
        68063 => X"14",  -- 20
        68064 => X"13",  -- 19
        68065 => X"19",  -- 25
        68066 => X"1D",  -- 29
        68067 => X"41",  -- 65
        68068 => X"60",  -- 96
        68069 => X"66",  -- 102
        68070 => X"75",  -- 117
        68071 => X"7B",  -- 123
        68072 => X"87",  -- 135
        68073 => X"91",  -- 145
        68074 => X"94",  -- 148
        68075 => X"8F",  -- 143
        68076 => X"8E",  -- 142
        68077 => X"92",  -- 146
        68078 => X"91",  -- 145
        68079 => X"88",  -- 136
        68080 => X"95",  -- 149
        68081 => X"81",  -- 129
        68082 => X"97",  -- 151
        68083 => X"94",  -- 148
        68084 => X"86",  -- 134
        68085 => X"92",  -- 146
        68086 => X"8C",  -- 140
        68087 => X"86",  -- 134
        68088 => X"7E",  -- 126
        68089 => X"7E",  -- 126
        68090 => X"74",  -- 116
        68091 => X"77",  -- 119
        68092 => X"8C",  -- 140
        68093 => X"93",  -- 147
        68094 => X"86",  -- 134
        68095 => X"7E",  -- 126
        68096 => X"84",  -- 132
        68097 => X"90",  -- 144
        68098 => X"90",  -- 144
        68099 => X"90",  -- 144
        68100 => X"9D",  -- 157
        68101 => X"98",  -- 152
        68102 => X"91",  -- 145
        68103 => X"96",  -- 150
        68104 => X"95",  -- 149
        68105 => X"8D",  -- 141
        68106 => X"82",  -- 130
        68107 => X"91",  -- 145
        68108 => X"96",  -- 150
        68109 => X"A6",  -- 166
        68110 => X"9D",  -- 157
        68111 => X"9B",  -- 155
        68112 => X"94",  -- 148
        68113 => X"8A",  -- 138
        68114 => X"A0",  -- 160
        68115 => X"A6",  -- 166
        68116 => X"A8",  -- 168
        68117 => X"BB",  -- 187
        68118 => X"B3",  -- 179
        68119 => X"9E",  -- 158
        68120 => X"89",  -- 137
        68121 => X"9C",  -- 156
        68122 => X"B8",  -- 184
        68123 => X"AE",  -- 174
        68124 => X"AC",  -- 172
        68125 => X"9E",  -- 158
        68126 => X"A6",  -- 166
        68127 => X"9F",  -- 159
        68128 => X"9F",  -- 159
        68129 => X"A2",  -- 162
        68130 => X"A8",  -- 168
        68131 => X"AA",  -- 170
        68132 => X"AE",  -- 174
        68133 => X"B1",  -- 177
        68134 => X"AE",  -- 174
        68135 => X"AA",  -- 170
        68136 => X"B4",  -- 180
        68137 => X"AF",  -- 175
        68138 => X"AB",  -- 171
        68139 => X"AC",  -- 172
        68140 => X"B0",  -- 176
        68141 => X"B0",  -- 176
        68142 => X"AD",  -- 173
        68143 => X"A8",  -- 168
        68144 => X"93",  -- 147
        68145 => X"96",  -- 150
        68146 => X"8D",  -- 141
        68147 => X"7E",  -- 126
        68148 => X"84",  -- 132
        68149 => X"89",  -- 137
        68150 => X"8D",  -- 141
        68151 => X"8F",  -- 143
        68152 => X"96",  -- 150
        68153 => X"81",  -- 129
        68154 => X"84",  -- 132
        68155 => X"84",  -- 132
        68156 => X"87",  -- 135
        68157 => X"9B",  -- 155
        68158 => X"9A",  -- 154
        68159 => X"8F",  -- 143
        68160 => X"72",  -- 114
        68161 => X"75",  -- 117
        68162 => X"77",  -- 119
        68163 => X"74",  -- 116
        68164 => X"70",  -- 112
        68165 => X"77",  -- 119
        68166 => X"7C",  -- 124
        68167 => X"74",  -- 116
        68168 => X"7B",  -- 123
        68169 => X"75",  -- 117
        68170 => X"6B",  -- 107
        68171 => X"67",  -- 103
        68172 => X"6F",  -- 111
        68173 => X"6F",  -- 111
        68174 => X"6F",  -- 111
        68175 => X"78",  -- 120
        68176 => X"6B",  -- 107
        68177 => X"5F",  -- 95
        68178 => X"70",  -- 112
        68179 => X"67",  -- 103
        68180 => X"61",  -- 97
        68181 => X"67",  -- 103
        68182 => X"5B",  -- 91
        68183 => X"6C",  -- 108
        68184 => X"65",  -- 101
        68185 => X"67",  -- 103
        68186 => X"72",  -- 114
        68187 => X"75",  -- 117
        68188 => X"63",  -- 99
        68189 => X"57",  -- 87
        68190 => X"73",  -- 115
        68191 => X"4F",  -- 79
        68192 => X"6B",  -- 107
        68193 => X"53",  -- 83
        68194 => X"90",  -- 144
        68195 => X"67",  -- 103
        68196 => X"58",  -- 88
        68197 => X"5A",  -- 90
        68198 => X"5D",  -- 93
        68199 => X"6A",  -- 106
        68200 => X"5A",  -- 90
        68201 => X"56",  -- 86
        68202 => X"56",  -- 86
        68203 => X"68",  -- 104
        68204 => X"93",  -- 147
        68205 => X"5D",  -- 93
        68206 => X"4C",  -- 76
        68207 => X"64",  -- 100
        68208 => X"94",  -- 148
        68209 => X"62",  -- 98
        68210 => X"4F",  -- 79
        68211 => X"6E",  -- 110
        68212 => X"50",  -- 80
        68213 => X"4E",  -- 78
        68214 => X"51",  -- 81
        68215 => X"4A",  -- 74
        68216 => X"48",  -- 72
        68217 => X"49",  -- 73
        68218 => X"57",  -- 87
        68219 => X"55",  -- 85
        68220 => X"52",  -- 82
        68221 => X"52",  -- 82
        68222 => X"49",  -- 73
        68223 => X"4B",  -- 75
        68224 => X"47",  -- 71
        68225 => X"44",  -- 68
        68226 => X"44",  -- 68
        68227 => X"47",  -- 71
        68228 => X"48",  -- 72
        68229 => X"44",  -- 68
        68230 => X"40",  -- 64
        68231 => X"3D",  -- 61
        68232 => X"35",  -- 53
        68233 => X"40",  -- 64
        68234 => X"3E",  -- 62
        68235 => X"41",  -- 65
        68236 => X"6B",  -- 107
        68237 => X"42",  -- 66
        68238 => X"27",  -- 39
        68239 => X"31",  -- 49
        68240 => X"2C",  -- 44
        68241 => X"2F",  -- 47
        68242 => X"2A",  -- 42
        68243 => X"33",  -- 51
        68244 => X"4A",  -- 74
        68245 => X"25",  -- 37
        68246 => X"2E",  -- 46
        68247 => X"31",  -- 49
        68248 => X"2A",  -- 42
        68249 => X"30",  -- 48
        68250 => X"39",  -- 57
        68251 => X"26",  -- 38
        68252 => X"3F",  -- 63
        68253 => X"2B",  -- 43
        68254 => X"1E",  -- 30
        68255 => X"2C",  -- 44
        68256 => X"2D",  -- 45
        68257 => X"2B",  -- 43
        68258 => X"59",  -- 89
        68259 => X"3E",  -- 62
        68260 => X"2F",  -- 47
        68261 => X"45",  -- 69
        68262 => X"30",  -- 48
        68263 => X"1D",  -- 29
        68264 => X"45",  -- 69
        68265 => X"25",  -- 37
        68266 => X"32",  -- 50
        68267 => X"3A",  -- 58
        68268 => X"27",  -- 39
        68269 => X"35",  -- 53
        68270 => X"4A",  -- 74
        68271 => X"54",  -- 84
        68272 => X"5A",  -- 90
        68273 => X"4D",  -- 77
        68274 => X"4D",  -- 77
        68275 => X"45",  -- 69
        68276 => X"39",  -- 57
        68277 => X"4A",  -- 74
        68278 => X"48",  -- 72
        68279 => X"21",  -- 33
        68280 => X"22",  -- 34
        68281 => X"1F",  -- 31
        68282 => X"17",  -- 23
        68283 => X"0F",  -- 15
        68284 => X"12",  -- 18
        68285 => X"1B",  -- 27
        68286 => X"1F",  -- 31
        68287 => X"1D",  -- 29
        68288 => X"20",  -- 32
        68289 => X"1D",  -- 29
        68290 => X"19",  -- 25
        68291 => X"35",  -- 53
        68292 => X"38",  -- 56
        68293 => X"3B",  -- 59
        68294 => X"49",  -- 73
        68295 => X"4B",  -- 75
        68296 => X"46",  -- 70
        68297 => X"2E",  -- 46
        68298 => X"25",  -- 37
        68299 => X"1F",  -- 31
        68300 => X"21",  -- 33
        68301 => X"5B",  -- 91
        68302 => X"5C",  -- 92
        68303 => X"0D",  -- 13
        68304 => X"12",  -- 18
        68305 => X"19",  -- 25
        68306 => X"2B",  -- 43
        68307 => X"58",  -- 88
        68308 => X"20",  -- 32
        68309 => X"3E",  -- 62
        68310 => X"49",  -- 73
        68311 => X"37",  -- 55
        68312 => X"34",  -- 52
        68313 => X"2A",  -- 42
        68314 => X"32",  -- 50
        68315 => X"36",  -- 54
        68316 => X"35",  -- 53
        68317 => X"30",  -- 48
        68318 => X"23",  -- 35
        68319 => X"2C",  -- 44
        68320 => X"3B",  -- 59
        68321 => X"3C",  -- 60
        68322 => X"75",  -- 117
        68323 => X"5C",  -- 92
        68324 => X"50",  -- 80
        68325 => X"53",  -- 83
        68326 => X"80",  -- 128
        68327 => X"4A",  -- 74
        68328 => X"4C",  -- 76
        68329 => X"4F",  -- 79
        68330 => X"4D",  -- 77
        68331 => X"4B",  -- 75
        68332 => X"50",  -- 80
        68333 => X"57",  -- 87
        68334 => X"58",  -- 88
        68335 => X"52",  -- 82
        68336 => X"44",  -- 68
        68337 => X"54",  -- 84
        68338 => X"5B",  -- 91
        68339 => X"5D",  -- 93
        68340 => X"5B",  -- 91
        68341 => X"55",  -- 85
        68342 => X"54",  -- 84
        68343 => X"5D",  -- 93
        68344 => X"5B",  -- 91
        68345 => X"63",  -- 99
        68346 => X"62",  -- 98
        68347 => X"5B",  -- 91
        68348 => X"5E",  -- 94
        68349 => X"6B",  -- 107
        68350 => X"6A",  -- 106
        68351 => X"5F",  -- 95
        68352 => X"5C",  -- 92
        68353 => X"5D",  -- 93
        68354 => X"62",  -- 98
        68355 => X"6B",  -- 107
        68356 => X"6F",  -- 111
        68357 => X"6D",  -- 109
        68358 => X"69",  -- 105
        68359 => X"67",  -- 103
        68360 => X"66",  -- 102
        68361 => X"5F",  -- 95
        68362 => X"62",  -- 98
        68363 => X"64",  -- 100
        68364 => X"5A",  -- 90
        68365 => X"52",  -- 82
        68366 => X"4F",  -- 79
        68367 => X"47",  -- 71
        68368 => X"3B",  -- 59
        68369 => X"36",  -- 54
        68370 => X"2E",  -- 46
        68371 => X"28",  -- 40
        68372 => X"23",  -- 35
        68373 => X"21",  -- 33
        68374 => X"22",  -- 34
        68375 => X"23",  -- 35
        68376 => X"24",  -- 36
        68377 => X"1D",  -- 29
        68378 => X"1A",  -- 26
        68379 => X"1D",  -- 29
        68380 => X"23",  -- 35
        68381 => X"26",  -- 38
        68382 => X"28",  -- 40
        68383 => X"2A",  -- 42
        68384 => X"33",  -- 51
        68385 => X"3E",  -- 62
        68386 => X"49",  -- 73
        68387 => X"76",  -- 118
        68388 => X"89",  -- 137
        68389 => X"7D",  -- 125
        68390 => X"88",  -- 136
        68391 => X"86",  -- 134
        68392 => X"97",  -- 151
        68393 => X"95",  -- 149
        68394 => X"93",  -- 147
        68395 => X"94",  -- 148
        68396 => X"9B",  -- 155
        68397 => X"9C",  -- 156
        68398 => X"91",  -- 145
        68399 => X"81",  -- 129
        68400 => X"8E",  -- 142
        68401 => X"84",  -- 132
        68402 => X"8F",  -- 143
        68403 => X"8E",  -- 142
        68404 => X"84",  -- 132
        68405 => X"8D",  -- 141
        68406 => X"92",  -- 146
        68407 => X"91",  -- 145
        68408 => X"91",  -- 145
        68409 => X"8B",  -- 139
        68410 => X"81",  -- 129
        68411 => X"89",  -- 137
        68412 => X"95",  -- 149
        68413 => X"89",  -- 137
        68414 => X"84",  -- 132
        68415 => X"9A",  -- 154
        68416 => X"94",  -- 148
        68417 => X"9A",  -- 154
        68418 => X"97",  -- 151
        68419 => X"96",  -- 150
        68420 => X"94",  -- 148
        68421 => X"8C",  -- 140
        68422 => X"81",  -- 129
        68423 => X"80",  -- 128
        68424 => X"93",  -- 147
        68425 => X"95",  -- 149
        68426 => X"97",  -- 151
        68427 => X"A3",  -- 163
        68428 => X"9D",  -- 157
        68429 => X"9C",  -- 156
        68430 => X"96",  -- 150
        68431 => X"9C",  -- 156
        68432 => X"8D",  -- 141
        68433 => X"92",  -- 146
        68434 => X"B5",  -- 181
        68435 => X"B3",  -- 179
        68436 => X"B8",  -- 184
        68437 => X"C4",  -- 196
        68438 => X"AC",  -- 172
        68439 => X"A0",  -- 160
        68440 => X"B4",  -- 180
        68441 => X"B2",  -- 178
        68442 => X"B5",  -- 181
        68443 => X"A7",  -- 167
        68444 => X"A3",  -- 163
        68445 => X"A5",  -- 165
        68446 => X"AB",  -- 171
        68447 => X"9D",  -- 157
        68448 => X"99",  -- 153
        68449 => X"A1",  -- 161
        68450 => X"A4",  -- 164
        68451 => X"A2",  -- 162
        68452 => X"A7",  -- 167
        68453 => X"AE",  -- 174
        68454 => X"AC",  -- 172
        68455 => X"A3",  -- 163
        68456 => X"A9",  -- 169
        68457 => X"A8",  -- 168
        68458 => X"AA",  -- 170
        68459 => X"B0",  -- 176
        68460 => X"B3",  -- 179
        68461 => X"A9",  -- 169
        68462 => X"93",  -- 147
        68463 => X"7F",  -- 127
        68464 => X"85",  -- 133
        68465 => X"8C",  -- 140
        68466 => X"90",  -- 144
        68467 => X"89",  -- 137
        68468 => X"96",  -- 150
        68469 => X"94",  -- 148
        68470 => X"99",  -- 153
        68471 => X"9B",  -- 155
        68472 => X"8D",  -- 141
        68473 => X"86",  -- 134
        68474 => X"91",  -- 145
        68475 => X"92",  -- 146
        68476 => X"96",  -- 150
        68477 => X"A1",  -- 161
        68478 => X"98",  -- 152
        68479 => X"91",  -- 145
        68480 => X"66",  -- 102
        68481 => X"73",  -- 115
        68482 => X"76",  -- 118
        68483 => X"6F",  -- 111
        68484 => X"70",  -- 112
        68485 => X"71",  -- 113
        68486 => X"71",  -- 113
        68487 => X"72",  -- 114
        68488 => X"6F",  -- 111
        68489 => X"70",  -- 112
        68490 => X"67",  -- 103
        68491 => X"63",  -- 99
        68492 => X"6C",  -- 108
        68493 => X"71",  -- 113
        68494 => X"6E",  -- 110
        68495 => X"6E",  -- 110
        68496 => X"56",  -- 86
        68497 => X"65",  -- 101
        68498 => X"6A",  -- 106
        68499 => X"62",  -- 98
        68500 => X"60",  -- 96
        68501 => X"54",  -- 84
        68502 => X"49",  -- 73
        68503 => X"57",  -- 87
        68504 => X"58",  -- 88
        68505 => X"56",  -- 86
        68506 => X"58",  -- 88
        68507 => X"5B",  -- 91
        68508 => X"55",  -- 85
        68509 => X"50",  -- 80
        68510 => X"6F",  -- 111
        68511 => X"56",  -- 86
        68512 => X"6F",  -- 111
        68513 => X"6D",  -- 109
        68514 => X"7C",  -- 124
        68515 => X"4E",  -- 78
        68516 => X"5B",  -- 91
        68517 => X"46",  -- 70
        68518 => X"5B",  -- 91
        68519 => X"58",  -- 88
        68520 => X"59",  -- 89
        68521 => X"4F",  -- 79
        68522 => X"46",  -- 70
        68523 => X"76",  -- 118
        68524 => X"66",  -- 102
        68525 => X"4C",  -- 76
        68526 => X"46",  -- 70
        68527 => X"74",  -- 116
        68528 => X"80",  -- 128
        68529 => X"4A",  -- 74
        68530 => X"56",  -- 86
        68531 => X"57",  -- 87
        68532 => X"3F",  -- 63
        68533 => X"4D",  -- 77
        68534 => X"48",  -- 72
        68535 => X"47",  -- 71
        68536 => X"46",  -- 70
        68537 => X"40",  -- 64
        68538 => X"51",  -- 81
        68539 => X"51",  -- 81
        68540 => X"4C",  -- 76
        68541 => X"4E",  -- 78
        68542 => X"40",  -- 64
        68543 => X"3F",  -- 63
        68544 => X"3B",  -- 59
        68545 => X"38",  -- 56
        68546 => X"37",  -- 55
        68547 => X"37",  -- 55
        68548 => X"36",  -- 54
        68549 => X"34",  -- 52
        68550 => X"35",  -- 53
        68551 => X"39",  -- 57
        68552 => X"2C",  -- 44
        68553 => X"3A",  -- 58
        68554 => X"32",  -- 50
        68555 => X"42",  -- 66
        68556 => X"4D",  -- 77
        68557 => X"32",  -- 50
        68558 => X"2C",  -- 44
        68559 => X"23",  -- 35
        68560 => X"26",  -- 38
        68561 => X"2C",  -- 44
        68562 => X"23",  -- 35
        68563 => X"23",  -- 35
        68564 => X"33",  -- 51
        68565 => X"26",  -- 38
        68566 => X"27",  -- 39
        68567 => X"2E",  -- 46
        68568 => X"20",  -- 32
        68569 => X"2B",  -- 43
        68570 => X"33",  -- 51
        68571 => X"25",  -- 37
        68572 => X"30",  -- 48
        68573 => X"2C",  -- 44
        68574 => X"1E",  -- 30
        68575 => X"25",  -- 37
        68576 => X"24",  -- 36
        68577 => X"31",  -- 49
        68578 => X"47",  -- 71
        68579 => X"2F",  -- 47
        68580 => X"27",  -- 39
        68581 => X"43",  -- 67
        68582 => X"23",  -- 35
        68583 => X"25",  -- 37
        68584 => X"2E",  -- 46
        68585 => X"1A",  -- 26
        68586 => X"2D",  -- 45
        68587 => X"32",  -- 50
        68588 => X"33",  -- 51
        68589 => X"3A",  -- 58
        68590 => X"44",  -- 68
        68591 => X"59",  -- 89
        68592 => X"4F",  -- 79
        68593 => X"47",  -- 71
        68594 => X"45",  -- 69
        68595 => X"3B",  -- 59
        68596 => X"2F",  -- 47
        68597 => X"3A",  -- 58
        68598 => X"3A",  -- 58
        68599 => X"1C",  -- 28
        68600 => X"12",  -- 18
        68601 => X"0F",  -- 15
        68602 => X"0A",  -- 10
        68603 => X"06",  -- 6
        68604 => X"05",  -- 5
        68605 => X"0A",  -- 10
        68606 => X"0F",  -- 15
        68607 => X"11",  -- 17
        68608 => X"10",  -- 16
        68609 => X"10",  -- 16
        68610 => X"0F",  -- 15
        68611 => X"1F",  -- 31
        68612 => X"20",  -- 32
        68613 => X"2D",  -- 45
        68614 => X"2E",  -- 46
        68615 => X"49",  -- 73
        68616 => X"27",  -- 39
        68617 => X"15",  -- 21
        68618 => X"0A",  -- 10
        68619 => X"08",  -- 8
        68620 => X"05",  -- 5
        68621 => X"31",  -- 49
        68622 => X"5E",  -- 94
        68623 => X"1C",  -- 28
        68624 => X"1E",  -- 30
        68625 => X"29",  -- 41
        68626 => X"33",  -- 51
        68627 => X"5C",  -- 92
        68628 => X"3D",  -- 61
        68629 => X"37",  -- 55
        68630 => X"44",  -- 68
        68631 => X"3D",  -- 61
        68632 => X"35",  -- 53
        68633 => X"2E",  -- 46
        68634 => X"3B",  -- 59
        68635 => X"3E",  -- 62
        68636 => X"38",  -- 56
        68637 => X"34",  -- 52
        68638 => X"39",  -- 57
        68639 => X"54",  -- 84
        68640 => X"3F",  -- 63
        68641 => X"44",  -- 68
        68642 => X"5A",  -- 90
        68643 => X"76",  -- 118
        68644 => X"4D",  -- 77
        68645 => X"4B",  -- 75
        68646 => X"68",  -- 104
        68647 => X"53",  -- 83
        68648 => X"4C",  -- 76
        68649 => X"50",  -- 80
        68650 => X"4E",  -- 78
        68651 => X"4C",  -- 76
        68652 => X"52",  -- 82
        68653 => X"5B",  -- 91
        68654 => X"5C",  -- 92
        68655 => X"56",  -- 86
        68656 => X"43",  -- 67
        68657 => X"55",  -- 85
        68658 => X"5F",  -- 95
        68659 => X"5F",  -- 95
        68660 => X"5A",  -- 90
        68661 => X"54",  -- 84
        68662 => X"56",  -- 86
        68663 => X"63",  -- 99
        68664 => X"64",  -- 100
        68665 => X"64",  -- 100
        68666 => X"61",  -- 97
        68667 => X"5F",  -- 95
        68668 => X"62",  -- 98
        68669 => X"67",  -- 103
        68670 => X"61",  -- 97
        68671 => X"56",  -- 86
        68672 => X"60",  -- 96
        68673 => X"5D",  -- 93
        68674 => X"61",  -- 97
        68675 => X"6C",  -- 108
        68676 => X"75",  -- 117
        68677 => X"75",  -- 117
        68678 => X"71",  -- 113
        68679 => X"6D",  -- 109
        68680 => X"63",  -- 99
        68681 => X"5B",  -- 91
        68682 => X"61",  -- 97
        68683 => X"69",  -- 105
        68684 => X"5D",  -- 93
        68685 => X"55",  -- 85
        68686 => X"4F",  -- 79
        68687 => X"43",  -- 67
        68688 => X"36",  -- 54
        68689 => X"35",  -- 53
        68690 => X"32",  -- 50
        68691 => X"30",  -- 48
        68692 => X"30",  -- 48
        68693 => X"30",  -- 48
        68694 => X"2E",  -- 46
        68695 => X"2D",  -- 45
        68696 => X"36",  -- 54
        68697 => X"31",  -- 49
        68698 => X"2F",  -- 47
        68699 => X"33",  -- 51
        68700 => X"37",  -- 55
        68701 => X"3A",  -- 58
        68702 => X"40",  -- 64
        68703 => X"46",  -- 70
        68704 => X"4E",  -- 78
        68705 => X"5F",  -- 95
        68706 => X"68",  -- 104
        68707 => X"8D",  -- 141
        68708 => X"91",  -- 145
        68709 => X"7F",  -- 127
        68710 => X"8C",  -- 140
        68711 => X"7F",  -- 127
        68712 => X"98",  -- 152
        68713 => X"8D",  -- 141
        68714 => X"86",  -- 134
        68715 => X"8B",  -- 139
        68716 => X"91",  -- 145
        68717 => X"8E",  -- 142
        68718 => X"84",  -- 132
        68719 => X"7B",  -- 123
        68720 => X"8C",  -- 140
        68721 => X"8F",  -- 143
        68722 => X"8A",  -- 138
        68723 => X"8D",  -- 141
        68724 => X"8B",  -- 139
        68725 => X"89",  -- 137
        68726 => X"93",  -- 147
        68727 => X"92",  -- 146
        68728 => X"89",  -- 137
        68729 => X"8B",  -- 139
        68730 => X"7B",  -- 123
        68731 => X"75",  -- 117
        68732 => X"80",  -- 128
        68733 => X"7C",  -- 124
        68734 => X"7E",  -- 126
        68735 => X"97",  -- 151
        68736 => X"99",  -- 153
        68737 => X"94",  -- 148
        68738 => X"96",  -- 150
        68739 => X"96",  -- 150
        68740 => X"91",  -- 145
        68741 => X"90",  -- 144
        68742 => X"92",  -- 146
        68743 => X"8D",  -- 141
        68744 => X"89",  -- 137
        68745 => X"8D",  -- 141
        68746 => X"91",  -- 145
        68747 => X"84",  -- 132
        68748 => X"7D",  -- 125
        68749 => X"77",  -- 119
        68750 => X"83",  -- 131
        68751 => X"8A",  -- 138
        68752 => X"A0",  -- 160
        68753 => X"A0",  -- 160
        68754 => X"9D",  -- 157
        68755 => X"9A",  -- 154
        68756 => X"AD",  -- 173
        68757 => X"B7",  -- 183
        68758 => X"B7",  -- 183
        68759 => X"C1",  -- 193
        68760 => X"AE",  -- 174
        68761 => X"A5",  -- 165
        68762 => X"A8",  -- 168
        68763 => X"B1",  -- 177
        68764 => X"AC",  -- 172
        68765 => X"B7",  -- 183
        68766 => X"B9",  -- 185
        68767 => X"B0",  -- 176
        68768 => X"AF",  -- 175
        68769 => X"A6",  -- 166
        68770 => X"A6",  -- 166
        68771 => X"AD",  -- 173
        68772 => X"AB",  -- 171
        68773 => X"A4",  -- 164
        68774 => X"A4",  -- 164
        68775 => X"AD",  -- 173
        68776 => X"A8",  -- 168
        68777 => X"99",  -- 153
        68778 => X"8F",  -- 143
        68779 => X"8F",  -- 143
        68780 => X"8D",  -- 141
        68781 => X"85",  -- 133
        68782 => X"80",  -- 128
        68783 => X"82",  -- 130
        68784 => X"85",  -- 133
        68785 => X"87",  -- 135
        68786 => X"8B",  -- 139
        68787 => X"83",  -- 131
        68788 => X"8F",  -- 143
        68789 => X"82",  -- 130
        68790 => X"87",  -- 135
        68791 => X"8D",  -- 141
        68792 => X"8B",  -- 139
        68793 => X"8C",  -- 140
        68794 => X"8C",  -- 140
        68795 => X"7F",  -- 127
        68796 => X"81",  -- 129
        68797 => X"8D",  -- 141
        68798 => X"91",  -- 145
        68799 => X"A2",  -- 162
        68800 => X"5F",  -- 95
        68801 => X"76",  -- 118
        68802 => X"77",  -- 119
        68803 => X"6B",  -- 107
        68804 => X"6A",  -- 106
        68805 => X"64",  -- 100
        68806 => X"5F",  -- 95
        68807 => X"66",  -- 102
        68808 => X"63",  -- 99
        68809 => X"6B",  -- 107
        68810 => X"65",  -- 101
        68811 => X"60",  -- 96
        68812 => X"6A",  -- 106
        68813 => X"71",  -- 113
        68814 => X"6D",  -- 109
        68815 => X"69",  -- 105
        68816 => X"5E",  -- 94
        68817 => X"6D",  -- 109
        68818 => X"61",  -- 97
        68819 => X"5F",  -- 95
        68820 => X"51",  -- 81
        68821 => X"45",  -- 69
        68822 => X"5B",  -- 91
        68823 => X"59",  -- 89
        68824 => X"61",  -- 97
        68825 => X"4F",  -- 79
        68826 => X"40",  -- 64
        68827 => X"43",  -- 67
        68828 => X"53",  -- 83
        68829 => X"5A",  -- 90
        68830 => X"7D",  -- 125
        68831 => X"69",  -- 105
        68832 => X"64",  -- 100
        68833 => X"8D",  -- 141
        68834 => X"4A",  -- 74
        68835 => X"4B",  -- 75
        68836 => X"4D",  -- 77
        68837 => X"47",  -- 71
        68838 => X"5A",  -- 90
        68839 => X"62",  -- 98
        68840 => X"5F",  -- 95
        68841 => X"56",  -- 86
        68842 => X"4B",  -- 75
        68843 => X"83",  -- 131
        68844 => X"39",  -- 57
        68845 => X"40",  -- 64
        68846 => X"43",  -- 67
        68847 => X"8E",  -- 142
        68848 => X"5A",  -- 90
        68849 => X"2B",  -- 43
        68850 => X"52",  -- 82
        68851 => X"34",  -- 52
        68852 => X"30",  -- 48
        68853 => X"4A",  -- 74
        68854 => X"43",  -- 67
        68855 => X"47",  -- 71
        68856 => X"3B",  -- 59
        68857 => X"30",  -- 48
        68858 => X"43",  -- 67
        68859 => X"46",  -- 70
        68860 => X"47",  -- 71
        68861 => X"4E",  -- 78
        68862 => X"3F",  -- 63
        68863 => X"3B",  -- 59
        68864 => X"35",  -- 53
        68865 => X"2A",  -- 42
        68866 => X"21",  -- 33
        68867 => X"21",  -- 33
        68868 => X"27",  -- 39
        68869 => X"2A",  -- 42
        68870 => X"2C",  -- 44
        68871 => X"2E",  -- 46
        68872 => X"34",  -- 52
        68873 => X"25",  -- 37
        68874 => X"1B",  -- 27
        68875 => X"59",  -- 89
        68876 => X"44",  -- 68
        68877 => X"21",  -- 33
        68878 => X"28",  -- 40
        68879 => X"27",  -- 39
        68880 => X"1D",  -- 29
        68881 => X"26",  -- 38
        68882 => X"1E",  -- 30
        68883 => X"19",  -- 25
        68884 => X"23",  -- 35
        68885 => X"24",  -- 36
        68886 => X"1D",  -- 29
        68887 => X"26",  -- 38
        68888 => X"1B",  -- 27
        68889 => X"23",  -- 35
        68890 => X"30",  -- 48
        68891 => X"28",  -- 40
        68892 => X"24",  -- 36
        68893 => X"31",  -- 49
        68894 => X"23",  -- 35
        68895 => X"14",  -- 20
        68896 => X"1B",  -- 27
        68897 => X"34",  -- 52
        68898 => X"2E",  -- 46
        68899 => X"24",  -- 36
        68900 => X"1C",  -- 28
        68901 => X"3D",  -- 61
        68902 => X"1C",  -- 28
        68903 => X"2E",  -- 46
        68904 => X"29",  -- 41
        68905 => X"17",  -- 23
        68906 => X"26",  -- 38
        68907 => X"1D",  -- 29
        68908 => X"35",  -- 53
        68909 => X"3A",  -- 58
        68910 => X"49",  -- 73
        68911 => X"64",  -- 100
        68912 => X"45",  -- 69
        68913 => X"41",  -- 65
        68914 => X"3A",  -- 58
        68915 => X"30",  -- 48
        68916 => X"2B",  -- 43
        68917 => X"2C",  -- 44
        68918 => X"27",  -- 39
        68919 => X"1D",  -- 29
        68920 => X"0B",  -- 11
        68921 => X"08",  -- 8
        68922 => X"05",  -- 5
        68923 => X"04",  -- 4
        68924 => X"03",  -- 3
        68925 => X"04",  -- 4
        68926 => X"0A",  -- 10
        68927 => X"11",  -- 17
        68928 => X"12",  -- 18
        68929 => X"0E",  -- 14
        68930 => X"18",  -- 24
        68931 => X"1A",  -- 26
        68932 => X"17",  -- 23
        68933 => X"26",  -- 38
        68934 => X"0C",  -- 12
        68935 => X"34",  -- 52
        68936 => X"15",  -- 21
        68937 => X"1E",  -- 30
        68938 => X"26",  -- 38
        68939 => X"2C",  -- 44
        68940 => X"24",  -- 36
        68941 => X"2E",  -- 46
        68942 => X"6A",  -- 106
        68943 => X"38",  -- 56
        68944 => X"33",  -- 51
        68945 => X"38",  -- 56
        68946 => X"2D",  -- 45
        68947 => X"56",  -- 86
        68948 => X"50",  -- 80
        68949 => X"3D",  -- 61
        68950 => X"33",  -- 51
        68951 => X"36",  -- 54
        68952 => X"3A",  -- 58
        68953 => X"3F",  -- 63
        68954 => X"47",  -- 71
        68955 => X"3D",  -- 61
        68956 => X"3F",  -- 63
        68957 => X"4B",  -- 75
        68958 => X"43",  -- 67
        68959 => X"3D",  -- 61
        68960 => X"48",  -- 72
        68961 => X"50",  -- 80
        68962 => X"4A",  -- 74
        68963 => X"78",  -- 120
        68964 => X"5F",  -- 95
        68965 => X"4B",  -- 75
        68966 => X"5F",  -- 95
        68967 => X"68",  -- 104
        68968 => X"3E",  -- 62
        68969 => X"4C",  -- 76
        68970 => X"57",  -- 87
        68971 => X"53",  -- 83
        68972 => X"52",  -- 82
        68973 => X"57",  -- 87
        68974 => X"5A",  -- 90
        68975 => X"59",  -- 89
        68976 => X"5E",  -- 94
        68977 => X"65",  -- 101
        68978 => X"64",  -- 100
        68979 => X"5D",  -- 93
        68980 => X"5D",  -- 93
        68981 => X"59",  -- 89
        68982 => X"58",  -- 88
        68983 => X"63",  -- 99
        68984 => X"5F",  -- 95
        68985 => X"5A",  -- 90
        68986 => X"5A",  -- 90
        68987 => X"61",  -- 97
        68988 => X"65",  -- 101
        68989 => X"62",  -- 98
        68990 => X"5A",  -- 90
        68991 => X"57",  -- 87
        68992 => X"62",  -- 98
        68993 => X"5D",  -- 93
        68994 => X"5F",  -- 95
        68995 => X"6B",  -- 107
        68996 => X"78",  -- 120
        68997 => X"7B",  -- 123
        68998 => X"77",  -- 119
        68999 => X"72",  -- 114
        69000 => X"64",  -- 100
        69001 => X"5B",  -- 91
        69002 => X"63",  -- 99
        69003 => X"6D",  -- 109
        69004 => X"62",  -- 98
        69005 => X"58",  -- 88
        69006 => X"52",  -- 82
        69007 => X"40",  -- 64
        69008 => X"45",  -- 69
        69009 => X"41",  -- 65
        69010 => X"3E",  -- 62
        69011 => X"3F",  -- 63
        69012 => X"40",  -- 64
        69013 => X"3C",  -- 60
        69014 => X"37",  -- 55
        69015 => X"32",  -- 50
        69016 => X"3F",  -- 63
        69017 => X"3C",  -- 60
        69018 => X"3F",  -- 63
        69019 => X"42",  -- 66
        69020 => X"43",  -- 67
        69021 => X"45",  -- 69
        69022 => X"4D",  -- 77
        69023 => X"56",  -- 86
        69024 => X"66",  -- 102
        69025 => X"7A",  -- 122
        69026 => X"7C",  -- 124
        69027 => X"92",  -- 146
        69028 => X"8D",  -- 141
        69029 => X"81",  -- 129
        69030 => X"94",  -- 148
        69031 => X"85",  -- 133
        69032 => X"7E",  -- 126
        69033 => X"7A",  -- 122
        69034 => X"7E",  -- 126
        69035 => X"88",  -- 136
        69036 => X"89",  -- 137
        69037 => X"80",  -- 128
        69038 => X"77",  -- 119
        69039 => X"75",  -- 117
        69040 => X"8E",  -- 142
        69041 => X"9A",  -- 154
        69042 => X"8B",  -- 139
        69043 => X"91",  -- 145
        69044 => X"93",  -- 147
        69045 => X"86",  -- 134
        69046 => X"8C",  -- 140
        69047 => X"85",  -- 133
        69048 => X"81",  -- 129
        69049 => X"9A",  -- 154
        69050 => X"8C",  -- 140
        69051 => X"77",  -- 119
        69052 => X"8C",  -- 140
        69053 => X"9C",  -- 156
        69054 => X"95",  -- 149
        69055 => X"91",  -- 145
        69056 => X"AD",  -- 173
        69057 => X"A0",  -- 160
        69058 => X"9F",  -- 159
        69059 => X"9B",  -- 155
        69060 => X"8E",  -- 142
        69061 => X"90",  -- 144
        69062 => X"97",  -- 151
        69063 => X"91",  -- 145
        69064 => X"8A",  -- 138
        69065 => X"8A",  -- 138
        69066 => X"88",  -- 136
        69067 => X"6C",  -- 108
        69068 => X"72",  -- 114
        69069 => X"7E",  -- 126
        69070 => X"9D",  -- 157
        69071 => X"A4",  -- 164
        69072 => X"A6",  -- 166
        69073 => X"AA",  -- 170
        69074 => X"8B",  -- 139
        69075 => X"9B",  -- 155
        69076 => X"B5",  -- 181
        69077 => X"A4",  -- 164
        69078 => X"9C",  -- 156
        69079 => X"99",  -- 153
        69080 => X"AA",  -- 170
        69081 => X"A3",  -- 163
        69082 => X"A8",  -- 168
        69083 => X"BF",  -- 191
        69084 => X"AC",  -- 172
        69085 => X"B0",  -- 176
        69086 => X"AF",  -- 175
        69087 => X"B0",  -- 176
        69088 => X"A0",  -- 160
        69089 => X"9C",  -- 156
        69090 => X"9B",  -- 155
        69091 => X"99",  -- 153
        69092 => X"94",  -- 148
        69093 => X"90",  -- 144
        69094 => X"96",  -- 150
        69095 => X"A2",  -- 162
        69096 => X"96",  -- 150
        69097 => X"87",  -- 135
        69098 => X"84",  -- 132
        69099 => X"91",  -- 145
        69100 => X"90",  -- 144
        69101 => X"83",  -- 131
        69102 => X"88",  -- 136
        69103 => X"9C",  -- 156
        69104 => X"8E",  -- 142
        69105 => X"87",  -- 135
        69106 => X"85",  -- 133
        69107 => X"79",  -- 121
        69108 => X"85",  -- 133
        69109 => X"78",  -- 120
        69110 => X"85",  -- 133
        69111 => X"93",  -- 147
        69112 => X"91",  -- 145
        69113 => X"91",  -- 145
        69114 => X"8C",  -- 140
        69115 => X"82",  -- 130
        69116 => X"90",  -- 144
        69117 => X"96",  -- 150
        69118 => X"86",  -- 134
        69119 => X"8B",  -- 139
        69120 => X"65",  -- 101
        69121 => X"58",  -- 88
        69122 => X"5E",  -- 94
        69123 => X"68",  -- 104
        69124 => X"5C",  -- 92
        69125 => X"4F",  -- 79
        69126 => X"5A",  -- 90
        69127 => X"6D",  -- 109
        69128 => X"70",  -- 112
        69129 => X"7B",  -- 123
        69130 => X"6F",  -- 111
        69131 => X"5C",  -- 92
        69132 => X"63",  -- 99
        69133 => X"71",  -- 113
        69134 => X"6B",  -- 107
        69135 => X"5C",  -- 92
        69136 => X"72",  -- 114
        69137 => X"6C",  -- 108
        69138 => X"61",  -- 97
        69139 => X"58",  -- 88
        69140 => X"53",  -- 83
        69141 => X"53",  -- 83
        69142 => X"56",  -- 86
        69143 => X"58",  -- 88
        69144 => X"50",  -- 80
        69145 => X"4A",  -- 74
        69146 => X"53",  -- 83
        69147 => X"4E",  -- 78
        69148 => X"59",  -- 89
        69149 => X"67",  -- 103
        69150 => X"82",  -- 130
        69151 => X"63",  -- 99
        69152 => X"6D",  -- 109
        69153 => X"66",  -- 102
        69154 => X"59",  -- 89
        69155 => X"4D",  -- 77
        69156 => X"4A",  -- 74
        69157 => X"4E",  -- 78
        69158 => X"53",  -- 83
        69159 => X"54",  -- 84
        69160 => X"6F",  -- 111
        69161 => X"52",  -- 82
        69162 => X"5F",  -- 95
        69163 => X"97",  -- 151
        69164 => X"38",  -- 56
        69165 => X"3D",  -- 61
        69166 => X"3F",  -- 63
        69167 => X"99",  -- 153
        69168 => X"44",  -- 68
        69169 => X"49",  -- 73
        69170 => X"56",  -- 86
        69171 => X"32",  -- 50
        69172 => X"3B",  -- 59
        69173 => X"2F",  -- 47
        69174 => X"44",  -- 68
        69175 => X"3B",  -- 59
        69176 => X"3D",  -- 61
        69177 => X"39",  -- 57
        69178 => X"4B",  -- 75
        69179 => X"47",  -- 71
        69180 => X"42",  -- 66
        69181 => X"45",  -- 69
        69182 => X"42",  -- 66
        69183 => X"56",  -- 86
        69184 => X"48",  -- 72
        69185 => X"2B",  -- 43
        69186 => X"1D",  -- 29
        69187 => X"20",  -- 32
        69188 => X"1F",  -- 31
        69189 => X"1E",  -- 30
        69190 => X"22",  -- 34
        69191 => X"23",  -- 35
        69192 => X"20",  -- 32
        69193 => X"20",  -- 32
        69194 => X"31",  -- 49
        69195 => X"54",  -- 84
        69196 => X"1F",  -- 31
        69197 => X"24",  -- 36
        69198 => X"21",  -- 33
        69199 => X"24",  -- 36
        69200 => X"1E",  -- 30
        69201 => X"1E",  -- 30
        69202 => X"22",  -- 34
        69203 => X"26",  -- 38
        69204 => X"25",  -- 37
        69205 => X"1F",  -- 31
        69206 => X"1D",  -- 29
        69207 => X"1D",  -- 29
        69208 => X"20",  -- 32
        69209 => X"26",  -- 38
        69210 => X"29",  -- 41
        69211 => X"27",  -- 39
        69212 => X"27",  -- 39
        69213 => X"28",  -- 40
        69214 => X"26",  -- 38
        69215 => X"21",  -- 33
        69216 => X"25",  -- 37
        69217 => X"2A",  -- 42
        69218 => X"2B",  -- 43
        69219 => X"15",  -- 21
        69220 => X"1D",  -- 29
        69221 => X"47",  -- 71
        69222 => X"25",  -- 37
        69223 => X"1C",  -- 28
        69224 => X"1F",  -- 31
        69225 => X"22",  -- 34
        69226 => X"1A",  -- 26
        69227 => X"14",  -- 20
        69228 => X"20",  -- 32
        69229 => X"33",  -- 51
        69230 => X"46",  -- 70
        69231 => X"57",  -- 87
        69232 => X"40",  -- 64
        69233 => X"43",  -- 67
        69234 => X"41",  -- 65
        69235 => X"32",  -- 50
        69236 => X"1F",  -- 31
        69237 => X"16",  -- 22
        69238 => X"1D",  -- 29
        69239 => X"27",  -- 39
        69240 => X"0E",  -- 14
        69241 => X"18",  -- 24
        69242 => X"1A",  -- 26
        69243 => X"11",  -- 17
        69244 => X"0B",  -- 11
        69245 => X"11",  -- 17
        69246 => X"1B",  -- 27
        69247 => X"1F",  -- 31
        69248 => X"25",  -- 37
        69249 => X"2A",  -- 42
        69250 => X"28",  -- 40
        69251 => X"22",  -- 34
        69252 => X"1C",  -- 28
        69253 => X"20",  -- 32
        69254 => X"22",  -- 34
        69255 => X"24",  -- 36
        69256 => X"30",  -- 48
        69257 => X"3F",  -- 63
        69258 => X"33",  -- 51
        69259 => X"38",  -- 56
        69260 => X"35",  -- 53
        69261 => X"3B",  -- 59
        69262 => X"62",  -- 98
        69263 => X"72",  -- 114
        69264 => X"34",  -- 52
        69265 => X"43",  -- 67
        69266 => X"3D",  -- 61
        69267 => X"46",  -- 70
        69268 => X"4D",  -- 77
        69269 => X"46",  -- 70
        69270 => X"3D",  -- 61
        69271 => X"32",  -- 50
        69272 => X"47",  -- 71
        69273 => X"43",  -- 67
        69274 => X"40",  -- 64
        69275 => X"42",  -- 66
        69276 => X"46",  -- 70
        69277 => X"48",  -- 72
        69278 => X"46",  -- 70
        69279 => X"43",  -- 67
        69280 => X"34",  -- 52
        69281 => X"4B",  -- 75
        69282 => X"44",  -- 68
        69283 => X"65",  -- 101
        69284 => X"81",  -- 129
        69285 => X"3A",  -- 58
        69286 => X"45",  -- 69
        69287 => X"77",  -- 119
        69288 => X"4C",  -- 76
        69289 => X"4A",  -- 74
        69290 => X"65",  -- 101
        69291 => X"55",  -- 85
        69292 => X"49",  -- 73
        69293 => X"51",  -- 81
        69294 => X"44",  -- 68
        69295 => X"59",  -- 89
        69296 => X"64",  -- 100
        69297 => X"60",  -- 96
        69298 => X"5B",  -- 91
        69299 => X"66",  -- 102
        69300 => X"5E",  -- 94
        69301 => X"49",  -- 73
        69302 => X"54",  -- 84
        69303 => X"60",  -- 96
        69304 => X"5D",  -- 93
        69305 => X"57",  -- 87
        69306 => X"57",  -- 87
        69307 => X"54",  -- 84
        69308 => X"5D",  -- 93
        69309 => X"61",  -- 97
        69310 => X"53",  -- 83
        69311 => X"5B",  -- 91
        69312 => X"62",  -- 98
        69313 => X"5F",  -- 95
        69314 => X"60",  -- 96
        69315 => X"65",  -- 101
        69316 => X"73",  -- 115
        69317 => X"7D",  -- 125
        69318 => X"79",  -- 121
        69319 => X"70",  -- 112
        69320 => X"67",  -- 103
        69321 => X"66",  -- 102
        69322 => X"64",  -- 100
        69323 => X"63",  -- 99
        69324 => X"62",  -- 98
        69325 => X"5B",  -- 91
        69326 => X"52",  -- 82
        69327 => X"4D",  -- 77
        69328 => X"4E",  -- 78
        69329 => X"4A",  -- 74
        69330 => X"4B",  -- 75
        69331 => X"50",  -- 80
        69332 => X"4D",  -- 77
        69333 => X"43",  -- 67
        69334 => X"42",  -- 66
        69335 => X"46",  -- 70
        69336 => X"45",  -- 69
        69337 => X"42",  -- 66
        69338 => X"42",  -- 66
        69339 => X"47",  -- 71
        69340 => X"4B",  -- 75
        69341 => X"51",  -- 81
        69342 => X"5F",  -- 95
        69343 => X"6C",  -- 108
        69344 => X"6E",  -- 110
        69345 => X"7C",  -- 124
        69346 => X"72",  -- 114
        69347 => X"7A",  -- 122
        69348 => X"7E",  -- 126
        69349 => X"68",  -- 104
        69350 => X"72",  -- 114
        69351 => X"95",  -- 149
        69352 => X"8A",  -- 138
        69353 => X"83",  -- 131
        69354 => X"81",  -- 129
        69355 => X"88",  -- 136
        69356 => X"8E",  -- 142
        69357 => X"8A",  -- 138
        69358 => X"83",  -- 131
        69359 => X"80",  -- 128
        69360 => X"7B",  -- 123
        69361 => X"74",  -- 116
        69362 => X"84",  -- 132
        69363 => X"89",  -- 137
        69364 => X"82",  -- 130
        69365 => X"84",  -- 132
        69366 => X"82",  -- 130
        69367 => X"87",  -- 135
        69368 => X"7D",  -- 125
        69369 => X"90",  -- 144
        69370 => X"94",  -- 148
        69371 => X"86",  -- 134
        69372 => X"90",  -- 144
        69373 => X"8D",  -- 141
        69374 => X"92",  -- 146
        69375 => X"77",  -- 119
        69376 => X"87",  -- 135
        69377 => X"81",  -- 129
        69378 => X"87",  -- 135
        69379 => X"96",  -- 150
        69380 => X"A0",  -- 160
        69381 => X"A2",  -- 162
        69382 => X"93",  -- 147
        69383 => X"7B",  -- 123
        69384 => X"89",  -- 137
        69385 => X"92",  -- 146
        69386 => X"77",  -- 119
        69387 => X"91",  -- 145
        69388 => X"93",  -- 147
        69389 => X"8B",  -- 139
        69390 => X"8A",  -- 138
        69391 => X"9A",  -- 154
        69392 => X"93",  -- 147
        69393 => X"9D",  -- 157
        69394 => X"A8",  -- 168
        69395 => X"A5",  -- 165
        69396 => X"B6",  -- 182
        69397 => X"8A",  -- 138
        69398 => X"A7",  -- 167
        69399 => X"AA",  -- 170
        69400 => X"A9",  -- 169
        69401 => X"B2",  -- 178
        69402 => X"A7",  -- 167
        69403 => X"A4",  -- 164
        69404 => X"90",  -- 144
        69405 => X"95",  -- 149
        69406 => X"83",  -- 131
        69407 => X"7C",  -- 124
        69408 => X"78",  -- 120
        69409 => X"79",  -- 121
        69410 => X"7D",  -- 125
        69411 => X"A0",  -- 160
        69412 => X"A8",  -- 168
        69413 => X"9B",  -- 155
        69414 => X"A6",  -- 166
        69415 => X"9E",  -- 158
        69416 => X"7B",  -- 123
        69417 => X"89",  -- 137
        69418 => X"7B",  -- 123
        69419 => X"87",  -- 135
        69420 => X"86",  -- 134
        69421 => X"93",  -- 147
        69422 => X"90",  -- 144
        69423 => X"93",  -- 147
        69424 => X"90",  -- 144
        69425 => X"8C",  -- 140
        69426 => X"81",  -- 129
        69427 => X"79",  -- 121
        69428 => X"86",  -- 134
        69429 => X"81",  -- 129
        69430 => X"91",  -- 145
        69431 => X"70",  -- 112
        69432 => X"82",  -- 130
        69433 => X"92",  -- 146
        69434 => X"7D",  -- 125
        69435 => X"98",  -- 152
        69436 => X"9A",  -- 154
        69437 => X"9D",  -- 157
        69438 => X"83",  -- 131
        69439 => X"A5",  -- 165
        69440 => X"5E",  -- 94
        69441 => X"58",  -- 88
        69442 => X"5F",  -- 95
        69443 => X"64",  -- 100
        69444 => X"59",  -- 89
        69445 => X"4C",  -- 76
        69446 => X"4F",  -- 79
        69447 => X"52",  -- 82
        69448 => X"69",  -- 105
        69449 => X"75",  -- 117
        69450 => X"6B",  -- 107
        69451 => X"55",  -- 85
        69452 => X"57",  -- 87
        69453 => X"65",  -- 101
        69454 => X"65",  -- 101
        69455 => X"60",  -- 96
        69456 => X"5E",  -- 94
        69457 => X"5F",  -- 95
        69458 => X"5E",  -- 94
        69459 => X"5C",  -- 92
        69460 => X"5A",  -- 90
        69461 => X"55",  -- 85
        69462 => X"53",  -- 83
        69463 => X"52",  -- 82
        69464 => X"50",  -- 80
        69465 => X"58",  -- 88
        69466 => X"5C",  -- 92
        69467 => X"63",  -- 99
        69468 => X"5A",  -- 90
        69469 => X"61",  -- 97
        69470 => X"73",  -- 115
        69471 => X"68",  -- 104
        69472 => X"75",  -- 117
        69473 => X"58",  -- 88
        69474 => X"47",  -- 71
        69475 => X"50",  -- 80
        69476 => X"52",  -- 82
        69477 => X"49",  -- 73
        69478 => X"4C",  -- 76
        69479 => X"5B",  -- 91
        69480 => X"67",  -- 103
        69481 => X"59",  -- 89
        69482 => X"7B",  -- 123
        69483 => X"6E",  -- 110
        69484 => X"39",  -- 57
        69485 => X"41",  -- 65
        69486 => X"53",  -- 83
        69487 => X"88",  -- 136
        69488 => X"3C",  -- 60
        69489 => X"48",  -- 72
        69490 => X"44",  -- 68
        69491 => X"2F",  -- 47
        69492 => X"2A",  -- 42
        69493 => X"37",  -- 55
        69494 => X"42",  -- 66
        69495 => X"3E",  -- 62
        69496 => X"3F",  -- 63
        69497 => X"39",  -- 57
        69498 => X"3D",  -- 61
        69499 => X"31",  -- 49
        69500 => X"35",  -- 53
        69501 => X"47",  -- 71
        69502 => X"43",  -- 67
        69503 => X"46",  -- 70
        69504 => X"40",  -- 64
        69505 => X"2C",  -- 44
        69506 => X"24",  -- 36
        69507 => X"25",  -- 37
        69508 => X"1E",  -- 30
        69509 => X"1C",  -- 28
        69510 => X"1D",  -- 29
        69511 => X"1A",  -- 26
        69512 => X"22",  -- 34
        69513 => X"1F",  -- 31
        69514 => X"32",  -- 50
        69515 => X"4F",  -- 79
        69516 => X"26",  -- 38
        69517 => X"25",  -- 37
        69518 => X"25",  -- 37
        69519 => X"25",  -- 37
        69520 => X"26",  -- 38
        69521 => X"21",  -- 33
        69522 => X"1F",  -- 31
        69523 => X"22",  -- 34
        69524 => X"24",  -- 36
        69525 => X"22",  -- 34
        69526 => X"1F",  -- 31
        69527 => X"1E",  -- 30
        69528 => X"22",  -- 34
        69529 => X"25",  -- 37
        69530 => X"22",  -- 34
        69531 => X"1C",  -- 28
        69532 => X"1A",  -- 26
        69533 => X"1D",  -- 29
        69534 => X"22",  -- 34
        69535 => X"24",  -- 36
        69536 => X"23",  -- 35
        69537 => X"1F",  -- 31
        69538 => X"20",  -- 32
        69539 => X"17",  -- 23
        69540 => X"1F",  -- 31
        69541 => X"3D",  -- 61
        69542 => X"1D",  -- 29
        69543 => X"1E",  -- 30
        69544 => X"1C",  -- 28
        69545 => X"20",  -- 32
        69546 => X"1A",  -- 26
        69547 => X"15",  -- 21
        69548 => X"1F",  -- 31
        69549 => X"2C",  -- 44
        69550 => X"36",  -- 54
        69551 => X"43",  -- 67
        69552 => X"4A",  -- 74
        69553 => X"42",  -- 66
        69554 => X"34",  -- 52
        69555 => X"23",  -- 35
        69556 => X"14",  -- 20
        69557 => X"10",  -- 16
        69558 => X"16",  -- 22
        69559 => X"1D",  -- 29
        69560 => X"1A",  -- 26
        69561 => X"1F",  -- 31
        69562 => X"21",  -- 33
        69563 => X"1D",  -- 29
        69564 => X"1D",  -- 29
        69565 => X"22",  -- 34
        69566 => X"2A",  -- 42
        69567 => X"2D",  -- 45
        69568 => X"35",  -- 53
        69569 => X"38",  -- 56
        69570 => X"38",  -- 56
        69571 => X"2F",  -- 47
        69572 => X"2C",  -- 44
        69573 => X"2F",  -- 47
        69574 => X"37",  -- 55
        69575 => X"3A",  -- 58
        69576 => X"3B",  -- 59
        69577 => X"34",  -- 52
        69578 => X"39",  -- 57
        69579 => X"41",  -- 65
        69580 => X"44",  -- 68
        69581 => X"3F",  -- 63
        69582 => X"54",  -- 84
        69583 => X"7F",  -- 127
        69584 => X"44",  -- 68
        69585 => X"3A",  -- 58
        69586 => X"3A",  -- 58
        69587 => X"4D",  -- 77
        69588 => X"53",  -- 83
        69589 => X"3B",  -- 59
        69590 => X"42",  -- 66
        69591 => X"47",  -- 71
        69592 => X"4F",  -- 79
        69593 => X"4C",  -- 76
        69594 => X"49",  -- 73
        69595 => X"48",  -- 72
        69596 => X"48",  -- 72
        69597 => X"47",  -- 71
        69598 => X"44",  -- 68
        69599 => X"40",  -- 64
        69600 => X"3C",  -- 60
        69601 => X"43",  -- 67
        69602 => X"43",  -- 67
        69603 => X"54",  -- 84
        69604 => X"6B",  -- 107
        69605 => X"52",  -- 82
        69606 => X"39",  -- 57
        69607 => X"61",  -- 97
        69608 => X"5B",  -- 91
        69609 => X"4E",  -- 78
        69610 => X"61",  -- 97
        69611 => X"5E",  -- 94
        69612 => X"5D",  -- 93
        69613 => X"5A",  -- 90
        69614 => X"39",  -- 57
        69615 => X"39",  -- 57
        69616 => X"55",  -- 85
        69617 => X"51",  -- 81
        69618 => X"4F",  -- 79
        69619 => X"5F",  -- 95
        69620 => X"56",  -- 86
        69621 => X"44",  -- 68
        69622 => X"63",  -- 99
        69623 => X"86",  -- 134
        69624 => X"68",  -- 104
        69625 => X"5C",  -- 92
        69626 => X"54",  -- 84
        69627 => X"4A",  -- 74
        69628 => X"54",  -- 84
        69629 => X"5B",  -- 91
        69630 => X"4F",  -- 79
        69631 => X"57",  -- 87
        69632 => X"60",  -- 96
        69633 => X"5E",  -- 94
        69634 => X"5D",  -- 93
        69635 => X"60",  -- 96
        69636 => X"6B",  -- 107
        69637 => X"74",  -- 116
        69638 => X"75",  -- 117
        69639 => X"70",  -- 112
        69640 => X"6A",  -- 106
        69641 => X"6B",  -- 107
        69642 => X"6A",  -- 106
        69643 => X"69",  -- 105
        69644 => X"66",  -- 102
        69645 => X"5E",  -- 94
        69646 => X"57",  -- 87
        69647 => X"52",  -- 82
        69648 => X"54",  -- 84
        69649 => X"51",  -- 81
        69650 => X"50",  -- 80
        69651 => X"54",  -- 84
        69652 => X"54",  -- 84
        69653 => X"52",  -- 82
        69654 => X"51",  -- 81
        69655 => X"52",  -- 82
        69656 => X"51",  -- 81
        69657 => X"50",  -- 80
        69658 => X"4D",  -- 77
        69659 => X"4E",  -- 78
        69660 => X"58",  -- 88
        69661 => X"67",  -- 103
        69662 => X"6E",  -- 110
        69663 => X"6E",  -- 110
        69664 => X"71",  -- 113
        69665 => X"8E",  -- 142
        69666 => X"80",  -- 128
        69667 => X"76",  -- 118
        69668 => X"7C",  -- 124
        69669 => X"7A",  -- 122
        69670 => X"7F",  -- 127
        69671 => X"84",  -- 132
        69672 => X"7A",  -- 122
        69673 => X"83",  -- 131
        69674 => X"8C",  -- 140
        69675 => X"8D",  -- 141
        69676 => X"83",  -- 131
        69677 => X"7F",  -- 127
        69678 => X"8A",  -- 138
        69679 => X"9B",  -- 155
        69680 => X"6F",  -- 111
        69681 => X"7C",  -- 124
        69682 => X"81",  -- 129
        69683 => X"8F",  -- 143
        69684 => X"7A",  -- 122
        69685 => X"78",  -- 120
        69686 => X"8C",  -- 140
        69687 => X"8B",  -- 139
        69688 => X"91",  -- 145
        69689 => X"96",  -- 150
        69690 => X"88",  -- 136
        69691 => X"7B",  -- 123
        69692 => X"93",  -- 147
        69693 => X"96",  -- 150
        69694 => X"9C",  -- 156
        69695 => X"88",  -- 136
        69696 => X"67",  -- 103
        69697 => X"77",  -- 119
        69698 => X"83",  -- 131
        69699 => X"83",  -- 131
        69700 => X"84",  -- 132
        69701 => X"8C",  -- 140
        69702 => X"94",  -- 148
        69703 => X"99",  -- 153
        69704 => X"9C",  -- 156
        69705 => X"9E",  -- 158
        69706 => X"89",  -- 137
        69707 => X"8C",  -- 140
        69708 => X"85",  -- 133
        69709 => X"6F",  -- 111
        69710 => X"85",  -- 133
        69711 => X"A6",  -- 166
        69712 => X"AD",  -- 173
        69713 => X"B3",  -- 179
        69714 => X"AD",  -- 173
        69715 => X"AA",  -- 170
        69716 => X"97",  -- 151
        69717 => X"A7",  -- 167
        69718 => X"A2",  -- 162
        69719 => X"C0",  -- 192
        69720 => X"C9",  -- 201
        69721 => X"BA",  -- 186
        69722 => X"A4",  -- 164
        69723 => X"A4",  -- 164
        69724 => X"8C",  -- 140
        69725 => X"84",  -- 132
        69726 => X"83",  -- 131
        69727 => X"99",  -- 153
        69728 => X"AB",  -- 171
        69729 => X"A6",  -- 166
        69730 => X"A5",  -- 165
        69731 => X"AF",  -- 175
        69732 => X"A9",  -- 169
        69733 => X"96",  -- 150
        69734 => X"8E",  -- 142
        69735 => X"83",  -- 131
        69736 => X"7E",  -- 126
        69737 => X"87",  -- 135
        69738 => X"81",  -- 129
        69739 => X"91",  -- 145
        69740 => X"90",  -- 144
        69741 => X"99",  -- 153
        69742 => X"95",  -- 149
        69743 => X"94",  -- 148
        69744 => X"90",  -- 144
        69745 => X"89",  -- 137
        69746 => X"71",  -- 113
        69747 => X"7E",  -- 126
        69748 => X"6A",  -- 106
        69749 => X"69",  -- 105
        69750 => X"71",  -- 113
        69751 => X"72",  -- 114
        69752 => X"60",  -- 96
        69753 => X"72",  -- 114
        69754 => X"74",  -- 116
        69755 => X"83",  -- 131
        69756 => X"76",  -- 118
        69757 => X"A3",  -- 163
        69758 => X"A4",  -- 164
        69759 => X"98",  -- 152
        69760 => X"58",  -- 88
        69761 => X"5B",  -- 91
        69762 => X"65",  -- 101
        69763 => X"69",  -- 105
        69764 => X"64",  -- 100
        69765 => X"63",  -- 99
        69766 => X"60",  -- 96
        69767 => X"56",  -- 86
        69768 => X"50",  -- 80
        69769 => X"68",  -- 104
        69770 => X"6B",  -- 107
        69771 => X"5C",  -- 92
        69772 => X"5C",  -- 92
        69773 => X"61",  -- 97
        69774 => X"61",  -- 97
        69775 => X"5F",  -- 95
        69776 => X"57",  -- 87
        69777 => X"5A",  -- 90
        69778 => X"5D",  -- 93
        69779 => X"5D",  -- 93
        69780 => X"5B",  -- 91
        69781 => X"57",  -- 87
        69782 => X"54",  -- 84
        69783 => X"52",  -- 82
        69784 => X"47",  -- 71
        69785 => X"52",  -- 82
        69786 => X"48",  -- 72
        69787 => X"59",  -- 89
        69788 => X"48",  -- 72
        69789 => X"4A",  -- 74
        69790 => X"54",  -- 84
        69791 => X"61",  -- 97
        69792 => X"6D",  -- 109
        69793 => X"4D",  -- 77
        69794 => X"3E",  -- 62
        69795 => X"4F",  -- 79
        69796 => X"5B",  -- 91
        69797 => X"53",  -- 83
        69798 => X"4D",  -- 77
        69799 => X"55",  -- 85
        69800 => X"58",  -- 88
        69801 => X"69",  -- 105
        69802 => X"92",  -- 146
        69803 => X"5E",  -- 94
        69804 => X"46",  -- 70
        69805 => X"4A",  -- 74
        69806 => X"5B",  -- 91
        69807 => X"66",  -- 102
        69808 => X"37",  -- 55
        69809 => X"45",  -- 69
        69810 => X"37",  -- 55
        69811 => X"37",  -- 55
        69812 => X"24",  -- 36
        69813 => X"40",  -- 64
        69814 => X"3A",  -- 58
        69815 => X"3A",  -- 58
        69816 => X"39",  -- 57
        69817 => X"3B",  -- 59
        69818 => X"3A",  -- 58
        69819 => X"28",  -- 40
        69820 => X"2D",  -- 45
        69821 => X"42",  -- 66
        69822 => X"3C",  -- 60
        69823 => X"30",  -- 48
        69824 => X"32",  -- 50
        69825 => X"2B",  -- 43
        69826 => X"2B",  -- 43
        69827 => X"2B",  -- 43
        69828 => X"25",  -- 37
        69829 => X"27",  -- 39
        69830 => X"29",  -- 41
        69831 => X"23",  -- 35
        69832 => X"20",  -- 32
        69833 => X"19",  -- 25
        69834 => X"30",  -- 48
        69835 => X"42",  -- 66
        69836 => X"2B",  -- 43
        69837 => X"23",  -- 35
        69838 => X"29",  -- 41
        69839 => X"24",  -- 36
        69840 => X"2A",  -- 42
        69841 => X"23",  -- 35
        69842 => X"20",  -- 32
        69843 => X"25",  -- 37
        69844 => X"2A",  -- 42
        69845 => X"28",  -- 40
        69846 => X"22",  -- 34
        69847 => X"1E",  -- 30
        69848 => X"22",  -- 34
        69849 => X"23",  -- 35
        69850 => X"21",  -- 33
        69851 => X"1B",  -- 27
        69852 => X"19",  -- 25
        69853 => X"1C",  -- 28
        69854 => X"21",  -- 33
        69855 => X"24",  -- 36
        69856 => X"25",  -- 37
        69857 => X"1A",  -- 26
        69858 => X"1A",  -- 26
        69859 => X"1E",  -- 30
        69860 => X"25",  -- 37
        69861 => X"34",  -- 52
        69862 => X"16",  -- 22
        69863 => X"20",  -- 32
        69864 => X"1C",  -- 28
        69865 => X"21",  -- 33
        69866 => X"1D",  -- 29
        69867 => X"1A",  -- 26
        69868 => X"21",  -- 33
        69869 => X"26",  -- 38
        69870 => X"27",  -- 39
        69871 => X"2C",  -- 44
        69872 => X"3B",  -- 59
        69873 => X"30",  -- 48
        69874 => X"20",  -- 32
        69875 => X"14",  -- 20
        69876 => X"13",  -- 19
        69877 => X"17",  -- 23
        69878 => X"1B",  -- 27
        69879 => X"1E",  -- 30
        69880 => X"25",  -- 37
        69881 => X"26",  -- 38
        69882 => X"27",  -- 39
        69883 => X"28",  -- 40
        69884 => X"2B",  -- 43
        69885 => X"32",  -- 50
        69886 => X"36",  -- 54
        69887 => X"37",  -- 55
        69888 => X"39",  -- 57
        69889 => X"3C",  -- 60
        69890 => X"38",  -- 56
        69891 => X"31",  -- 49
        69892 => X"2D",  -- 45
        69893 => X"33",  -- 51
        69894 => X"3D",  -- 61
        69895 => X"45",  -- 69
        69896 => X"45",  -- 69
        69897 => X"38",  -- 56
        69898 => X"43",  -- 67
        69899 => X"43",  -- 67
        69900 => X"45",  -- 69
        69901 => X"41",  -- 65
        69902 => X"3D",  -- 61
        69903 => X"73",  -- 115
        69904 => X"51",  -- 81
        69905 => X"3B",  -- 59
        69906 => X"42",  -- 66
        69907 => X"51",  -- 81
        69908 => X"59",  -- 89
        69909 => X"35",  -- 53
        69910 => X"44",  -- 68
        69911 => X"48",  -- 72
        69912 => X"47",  -- 71
        69913 => X"47",  -- 71
        69914 => X"48",  -- 72
        69915 => X"48",  -- 72
        69916 => X"48",  -- 72
        69917 => X"48",  -- 72
        69918 => X"47",  -- 71
        69919 => X"47",  -- 71
        69920 => X"47",  -- 71
        69921 => X"40",  -- 64
        69922 => X"4C",  -- 76
        69923 => X"49",  -- 73
        69924 => X"4E",  -- 78
        69925 => X"61",  -- 97
        69926 => X"2F",  -- 47
        69927 => X"49",  -- 73
        69928 => X"76",  -- 118
        69929 => X"55",  -- 85
        69930 => X"4E",  -- 78
        69931 => X"48",  -- 72
        69932 => X"50",  -- 80
        69933 => X"58",  -- 88
        69934 => X"47",  -- 71
        69935 => X"51",  -- 81
        69936 => X"58",  -- 88
        69937 => X"53",  -- 83
        69938 => X"54",  -- 84
        69939 => X"6A",  -- 106
        69940 => X"63",  -- 99
        69941 => X"4F",  -- 79
        69942 => X"67",  -- 103
        69943 => X"88",  -- 136
        69944 => X"6D",  -- 109
        69945 => X"5E",  -- 94
        69946 => X"52",  -- 82
        69947 => X"49",  -- 73
        69948 => X"57",  -- 87
        69949 => X"63",  -- 99
        69950 => X"59",  -- 89
        69951 => X"5D",  -- 93
        69952 => X"5A",  -- 90
        69953 => X"59",  -- 89
        69954 => X"57",  -- 87
        69955 => X"57",  -- 87
        69956 => X"5F",  -- 95
        69957 => X"68",  -- 104
        69958 => X"6E",  -- 110
        69959 => X"6E",  -- 110
        69960 => X"6C",  -- 108
        69961 => X"6F",  -- 111
        69962 => X"71",  -- 113
        69963 => X"6D",  -- 109
        69964 => X"67",  -- 103
        69965 => X"5E",  -- 94
        69966 => X"59",  -- 89
        69967 => X"57",  -- 87
        69968 => X"56",  -- 86
        69969 => X"57",  -- 87
        69970 => X"55",  -- 85
        69971 => X"56",  -- 86
        69972 => X"5A",  -- 90
        69973 => X"5F",  -- 95
        69974 => X"5F",  -- 95
        69975 => X"5C",  -- 92
        69976 => X"5D",  -- 93
        69977 => X"65",  -- 101
        69978 => X"63",  -- 99
        69979 => X"5C",  -- 92
        69980 => X"63",  -- 99
        69981 => X"73",  -- 115
        69982 => X"77",  -- 119
        69983 => X"6F",  -- 111
        69984 => X"74",  -- 116
        69985 => X"8D",  -- 141
        69986 => X"7E",  -- 126
        69987 => X"72",  -- 114
        69988 => X"80",  -- 128
        69989 => X"88",  -- 136
        69990 => X"89",  -- 137
        69991 => X"7F",  -- 127
        69992 => X"89",  -- 137
        69993 => X"85",  -- 133
        69994 => X"7F",  -- 127
        69995 => X"7A",  -- 122
        69996 => X"74",  -- 116
        69997 => X"6C",  -- 108
        69998 => X"67",  -- 103
        69999 => X"68",  -- 104
        70000 => X"7D",  -- 125
        70001 => X"8A",  -- 138
        70002 => X"6E",  -- 110
        70003 => X"79",  -- 121
        70004 => X"5D",  -- 93
        70005 => X"65",  -- 101
        70006 => X"8A",  -- 138
        70007 => X"81",  -- 129
        70008 => X"7F",  -- 127
        70009 => X"80",  -- 128
        70010 => X"6E",  -- 110
        70011 => X"6A",  -- 106
        70012 => X"8C",  -- 140
        70013 => X"8D",  -- 141
        70014 => X"92",  -- 146
        70015 => X"88",  -- 136
        70016 => X"74",  -- 116
        70017 => X"7A",  -- 122
        70018 => X"7E",  -- 126
        70019 => X"8A",  -- 138
        70020 => X"96",  -- 150
        70021 => X"8C",  -- 140
        70022 => X"8C",  -- 140
        70023 => X"A2",  -- 162
        70024 => X"8D",  -- 141
        70025 => X"91",  -- 145
        70026 => X"81",  -- 129
        70027 => X"8A",  -- 138
        70028 => X"77",  -- 119
        70029 => X"66",  -- 102
        70030 => X"72",  -- 114
        70031 => X"94",  -- 148
        70032 => X"B0",  -- 176
        70033 => X"AB",  -- 171
        70034 => X"AC",  -- 172
        70035 => X"A2",  -- 162
        70036 => X"8C",  -- 140
        70037 => X"B3",  -- 179
        70038 => X"84",  -- 132
        70039 => X"9E",  -- 158
        70040 => X"BB",  -- 187
        70041 => X"A2",  -- 162
        70042 => X"81",  -- 129
        70043 => X"83",  -- 131
        70044 => X"92",  -- 146
        70045 => X"AD",  -- 173
        70046 => X"AA",  -- 170
        70047 => X"A3",  -- 163
        70048 => X"97",  -- 151
        70049 => X"A4",  -- 164
        70050 => X"B4",  -- 180
        70051 => X"A3",  -- 163
        70052 => X"85",  -- 133
        70053 => X"77",  -- 119
        70054 => X"73",  -- 115
        70055 => X"80",  -- 128
        70056 => X"78",  -- 120
        70057 => X"91",  -- 145
        70058 => X"93",  -- 147
        70059 => X"87",  -- 135
        70060 => X"81",  -- 129
        70061 => X"A2",  -- 162
        70062 => X"9A",  -- 154
        70063 => X"7A",  -- 122
        70064 => X"55",  -- 85
        70065 => X"4A",  -- 74
        70066 => X"46",  -- 70
        70067 => X"6E",  -- 110
        70068 => X"64",  -- 100
        70069 => X"5E",  -- 94
        70070 => X"66",  -- 102
        70071 => X"76",  -- 118
        70072 => X"6C",  -- 108
        70073 => X"66",  -- 102
        70074 => X"5F",  -- 95
        70075 => X"71",  -- 113
        70076 => X"60",  -- 96
        70077 => X"76",  -- 118
        70078 => X"78",  -- 120
        70079 => X"7B",  -- 123
        70080 => X"50",  -- 80
        70081 => X"57",  -- 87
        70082 => X"5F",  -- 95
        70083 => X"5F",  -- 95
        70084 => X"61",  -- 97
        70085 => X"6E",  -- 110
        70086 => X"6D",  -- 109
        70087 => X"5B",  -- 91
        70088 => X"51",  -- 81
        70089 => X"68",  -- 104
        70090 => X"6C",  -- 108
        70091 => X"60",  -- 96
        70092 => X"5C",  -- 92
        70093 => X"5D",  -- 93
        70094 => X"5B",  -- 91
        70095 => X"5A",  -- 90
        70096 => X"5B",  -- 91
        70097 => X"5A",  -- 90
        70098 => X"58",  -- 88
        70099 => X"53",  -- 83
        70100 => X"51",  -- 81
        70101 => X"50",  -- 80
        70102 => X"53",  -- 83
        70103 => X"56",  -- 86
        70104 => X"52",  -- 82
        70105 => X"51",  -- 81
        70106 => X"3F",  -- 63
        70107 => X"4B",  -- 75
        70108 => X"47",  -- 71
        70109 => X"45",  -- 69
        70110 => X"55",  -- 85
        70111 => X"6D",  -- 109
        70112 => X"52",  -- 82
        70113 => X"4C",  -- 76
        70114 => X"46",  -- 70
        70115 => X"4A",  -- 74
        70116 => X"59",  -- 89
        70117 => X"63",  -- 99
        70118 => X"57",  -- 87
        70119 => X"44",  -- 68
        70120 => X"4A",  -- 74
        70121 => X"79",  -- 121
        70122 => X"84",  -- 132
        70123 => X"5A",  -- 90
        70124 => X"47",  -- 71
        70125 => X"4C",  -- 76
        70126 => X"64",  -- 100
        70127 => X"55",  -- 85
        70128 => X"33",  -- 51
        70129 => X"3A",  -- 58
        70130 => X"30",  -- 48
        70131 => X"40",  -- 64
        70132 => X"2E",  -- 46
        70133 => X"3B",  -- 59
        70134 => X"28",  -- 40
        70135 => X"29",  -- 41
        70136 => X"22",  -- 34
        70137 => X"31",  -- 49
        70138 => X"3B",  -- 59
        70139 => X"34",  -- 52
        70140 => X"34",  -- 52
        70141 => X"3D",  -- 61
        70142 => X"37",  -- 55
        70143 => X"2A",  -- 42
        70144 => X"2A",  -- 42
        70145 => X"28",  -- 40
        70146 => X"2B",  -- 43
        70147 => X"2A",  -- 42
        70148 => X"27",  -- 39
        70149 => X"30",  -- 48
        70150 => X"34",  -- 52
        70151 => X"2A",  -- 42
        70152 => X"1D",  -- 29
        70153 => X"13",  -- 19
        70154 => X"2C",  -- 44
        70155 => X"33",  -- 51
        70156 => X"2E",  -- 46
        70157 => X"20",  -- 32
        70158 => X"2A",  -- 42
        70159 => X"22",  -- 34
        70160 => X"24",  -- 36
        70161 => X"21",  -- 33
        70162 => X"22",  -- 34
        70163 => X"2A",  -- 42
        70164 => X"2E",  -- 46
        70165 => X"2A",  -- 42
        70166 => X"23",  -- 35
        70167 => X"1F",  -- 31
        70168 => X"1F",  -- 31
        70169 => X"1F",  -- 31
        70170 => X"1F",  -- 31
        70171 => X"20",  -- 32
        70172 => X"21",  -- 33
        70173 => X"21",  -- 33
        70174 => X"1E",  -- 30
        70175 => X"1A",  -- 26
        70176 => X"20",  -- 32
        70177 => X"1A",  -- 26
        70178 => X"18",  -- 24
        70179 => X"20",  -- 32
        70180 => X"23",  -- 35
        70181 => X"2D",  -- 45
        70182 => X"15",  -- 21
        70183 => X"1D",  -- 29
        70184 => X"1C",  -- 28
        70185 => X"22",  -- 34
        70186 => X"1E",  -- 30
        70187 => X"1B",  -- 27
        70188 => X"21",  -- 33
        70189 => X"21",  -- 33
        70190 => X"1B",  -- 27
        70191 => X"1A",  -- 26
        70192 => X"1F",  -- 31
        70193 => X"19",  -- 25
        70194 => X"15",  -- 21
        70195 => X"17",  -- 23
        70196 => X"20",  -- 32
        70197 => X"26",  -- 38
        70198 => X"26",  -- 38
        70199 => X"22",  -- 34
        70200 => X"2B",  -- 43
        70201 => X"2B",  -- 43
        70202 => X"2D",  -- 45
        70203 => X"30",  -- 48
        70204 => X"32",  -- 50
        70205 => X"33",  -- 51
        70206 => X"35",  -- 53
        70207 => X"39",  -- 57
        70208 => X"3B",  -- 59
        70209 => X"36",  -- 54
        70210 => X"2F",  -- 47
        70211 => X"28",  -- 40
        70212 => X"28",  -- 40
        70213 => X"2E",  -- 46
        70214 => X"38",  -- 56
        70215 => X"3E",  -- 62
        70216 => X"47",  -- 71
        70217 => X"47",  -- 71
        70218 => X"45",  -- 69
        70219 => X"3B",  -- 59
        70220 => X"40",  -- 64
        70221 => X"40",  -- 64
        70222 => X"3A",  -- 58
        70223 => X"59",  -- 89
        70224 => X"4F",  -- 79
        70225 => X"3D",  -- 61
        70226 => X"4A",  -- 74
        70227 => X"4E",  -- 78
        70228 => X"5C",  -- 92
        70229 => X"3A",  -- 58
        70230 => X"4A",  -- 74
        70231 => X"3B",  -- 59
        70232 => X"3A",  -- 58
        70233 => X"3D",  -- 61
        70234 => X"41",  -- 65
        70235 => X"43",  -- 67
        70236 => X"43",  -- 67
        70237 => X"45",  -- 69
        70238 => X"47",  -- 71
        70239 => X"49",  -- 73
        70240 => X"4A",  -- 74
        70241 => X"41",  -- 65
        70242 => X"57",  -- 87
        70243 => X"48",  -- 72
        70244 => X"46",  -- 70
        70245 => X"60",  -- 96
        70246 => X"3C",  -- 60
        70247 => X"4F",  -- 79
        70248 => X"5A",  -- 90
        70249 => X"44",  -- 68
        70250 => X"4A",  -- 74
        70251 => X"52",  -- 82
        70252 => X"5A",  -- 90
        70253 => X"5B",  -- 91
        70254 => X"4F",  -- 79
        70255 => X"5B",  -- 91
        70256 => X"57",  -- 87
        70257 => X"4B",  -- 75
        70258 => X"43",  -- 67
        70259 => X"56",  -- 86
        70260 => X"58",  -- 88
        70261 => X"49",  -- 73
        70262 => X"50",  -- 80
        70263 => X"59",  -- 89
        70264 => X"62",  -- 98
        70265 => X"54",  -- 84
        70266 => X"4B",  -- 75
        70267 => X"44",  -- 68
        70268 => X"55",  -- 85
        70269 => X"62",  -- 98
        70270 => X"54",  -- 84
        70271 => X"53",  -- 83
        70272 => X"59",  -- 89
        70273 => X"5A",  -- 90
        70274 => X"5A",  -- 90
        70275 => X"58",  -- 88
        70276 => X"5C",  -- 92
        70277 => X"65",  -- 101
        70278 => X"6D",  -- 109
        70279 => X"6F",  -- 111
        70280 => X"6E",  -- 110
        70281 => X"72",  -- 114
        70282 => X"73",  -- 115
        70283 => X"6F",  -- 111
        70284 => X"64",  -- 100
        70285 => X"5C",  -- 92
        70286 => X"59",  -- 89
        70287 => X"59",  -- 89
        70288 => X"57",  -- 87
        70289 => X"5B",  -- 91
        70290 => X"5B",  -- 91
        70291 => X"55",  -- 85
        70292 => X"56",  -- 86
        70293 => X"5D",  -- 93
        70294 => X"5F",  -- 95
        70295 => X"5C",  -- 92
        70296 => X"5E",  -- 94
        70297 => X"6E",  -- 110
        70298 => X"74",  -- 116
        70299 => X"6C",  -- 108
        70300 => X"66",  -- 102
        70301 => X"6B",  -- 107
        70302 => X"72",  -- 114
        70303 => X"74",  -- 116
        70304 => X"82",  -- 130
        70305 => X"82",  -- 130
        70306 => X"6F",  -- 111
        70307 => X"77",  -- 119
        70308 => X"88",  -- 136
        70309 => X"83",  -- 131
        70310 => X"81",  -- 129
        70311 => X"7E",  -- 126
        70312 => X"83",  -- 131
        70313 => X"74",  -- 116
        70314 => X"6C",  -- 108
        70315 => X"71",  -- 113
        70316 => X"7C",  -- 124
        70317 => X"7E",  -- 126
        70318 => X"6E",  -- 110
        70319 => X"5E",  -- 94
        70320 => X"79",  -- 121
        70321 => X"82",  -- 130
        70322 => X"69",  -- 105
        70323 => X"78",  -- 120
        70324 => X"68",  -- 104
        70325 => X"74",  -- 116
        70326 => X"77",  -- 119
        70327 => X"58",  -- 88
        70328 => X"6B",  -- 107
        70329 => X"72",  -- 114
        70330 => X"6B",  -- 107
        70331 => X"71",  -- 113
        70332 => X"93",  -- 147
        70333 => X"89",  -- 137
        70334 => X"8A",  -- 138
        70335 => X"87",  -- 135
        70336 => X"8D",  -- 141
        70337 => X"8C",  -- 140
        70338 => X"74",  -- 116
        70339 => X"69",  -- 105
        70340 => X"76",  -- 118
        70341 => X"79",  -- 121
        70342 => X"82",  -- 130
        70343 => X"A1",  -- 161
        70344 => X"8E",  -- 142
        70345 => X"91",  -- 145
        70346 => X"7F",  -- 127
        70347 => X"99",  -- 153
        70348 => X"87",  -- 135
        70349 => X"8F",  -- 143
        70350 => X"80",  -- 128
        70351 => X"8E",  -- 142
        70352 => X"9C",  -- 156
        70353 => X"93",  -- 147
        70354 => X"AA",  -- 170
        70355 => X"8D",  -- 141
        70356 => X"8B",  -- 139
        70357 => X"8B",  -- 139
        70358 => X"6D",  -- 109
        70359 => X"7C",  -- 124
        70360 => X"9A",  -- 154
        70361 => X"9C",  -- 156
        70362 => X"93",  -- 147
        70363 => X"8C",  -- 140
        70364 => X"92",  -- 146
        70365 => X"A6",  -- 166
        70366 => X"A9",  -- 169
        70367 => X"A2",  -- 162
        70368 => X"93",  -- 147
        70369 => X"8C",  -- 140
        70370 => X"8F",  -- 143
        70371 => X"83",  -- 131
        70372 => X"86",  -- 134
        70373 => X"8D",  -- 141
        70374 => X"78",  -- 120
        70375 => X"7B",  -- 123
        70376 => X"79",  -- 121
        70377 => X"85",  -- 133
        70378 => X"85",  -- 133
        70379 => X"6A",  -- 106
        70380 => X"61",  -- 97
        70381 => X"7A",  -- 122
        70382 => X"6F",  -- 111
        70383 => X"4A",  -- 74
        70384 => X"54",  -- 84
        70385 => X"33",  -- 51
        70386 => X"36",  -- 54
        70387 => X"47",  -- 71
        70388 => X"57",  -- 87
        70389 => X"42",  -- 66
        70390 => X"53",  -- 83
        70391 => X"5C",  -- 92
        70392 => X"65",  -- 101
        70393 => X"60",  -- 96
        70394 => X"43",  -- 67
        70395 => X"54",  -- 84
        70396 => X"5F",  -- 95
        70397 => X"5A",  -- 90
        70398 => X"54",  -- 84
        70399 => X"84",  -- 132
        70400 => X"59",  -- 89
        70401 => X"5C",  -- 92
        70402 => X"5D",  -- 93
        70403 => X"55",  -- 85
        70404 => X"55",  -- 85
        70405 => X"67",  -- 103
        70406 => X"6D",  -- 109
        70407 => X"5D",  -- 93
        70408 => X"69",  -- 105
        70409 => X"70",  -- 112
        70410 => X"65",  -- 101
        70411 => X"54",  -- 84
        70412 => X"51",  -- 81
        70413 => X"54",  -- 84
        70414 => X"55",  -- 85
        70415 => X"58",  -- 88
        70416 => X"58",  -- 88
        70417 => X"56",  -- 86
        70418 => X"50",  -- 80
        70419 => X"4A",  -- 74
        70420 => X"47",  -- 71
        70421 => X"48",  -- 72
        70422 => X"50",  -- 80
        70423 => X"56",  -- 86
        70424 => X"5A",  -- 90
        70425 => X"54",  -- 84
        70426 => X"4C",  -- 76
        70427 => X"49",  -- 73
        70428 => X"50",  -- 80
        70429 => X"43",  -- 67
        70430 => X"63",  -- 99
        70431 => X"7E",  -- 126
        70432 => X"42",  -- 66
        70433 => X"4A",  -- 74
        70434 => X"47",  -- 71
        70435 => X"41",  -- 65
        70436 => X"50",  -- 80
        70437 => X"62",  -- 98
        70438 => X"58",  -- 88
        70439 => X"3F",  -- 63
        70440 => X"47",  -- 71
        70441 => X"87",  -- 135
        70442 => X"6F",  -- 111
        70443 => X"43",  -- 67
        70444 => X"3E",  -- 62
        70445 => X"46",  -- 70
        70446 => X"82",  -- 130
        70447 => X"54",  -- 84
        70448 => X"34",  -- 52
        70449 => X"2B",  -- 43
        70450 => X"2B",  -- 43
        70451 => X"3D",  -- 61
        70452 => X"38",  -- 56
        70453 => X"29",  -- 41
        70454 => X"1A",  -- 26
        70455 => X"1D",  -- 29
        70456 => X"11",  -- 17
        70457 => X"1D",  -- 29
        70458 => X"2A",  -- 42
        70459 => X"39",  -- 57
        70460 => X"3E",  -- 62
        70461 => X"39",  -- 57
        70462 => X"34",  -- 52
        70463 => X"2B",  -- 43
        70464 => X"29",  -- 41
        70465 => X"24",  -- 36
        70466 => X"21",  -- 33
        70467 => X"1E",  -- 30
        70468 => X"1F",  -- 31
        70469 => X"2B",  -- 43
        70470 => X"2F",  -- 47
        70471 => X"23",  -- 35
        70472 => X"23",  -- 35
        70473 => X"19",  -- 25
        70474 => X"2F",  -- 47
        70475 => X"2E",  -- 46
        70476 => X"30",  -- 48
        70477 => X"1F",  -- 31
        70478 => X"28",  -- 40
        70479 => X"1F",  -- 31
        70480 => X"1E",  -- 30
        70481 => X"1D",  -- 29
        70482 => X"1F",  -- 31
        70483 => X"25",  -- 37
        70484 => X"26",  -- 38
        70485 => X"24",  -- 36
        70486 => X"23",  -- 35
        70487 => X"24",  -- 36
        70488 => X"22",  -- 34
        70489 => X"1D",  -- 29
        70490 => X"1B",  -- 27
        70491 => X"1F",  -- 31
        70492 => X"22",  -- 34
        70493 => X"1F",  -- 31
        70494 => X"16",  -- 22
        70495 => X"0D",  -- 13
        70496 => X"14",  -- 20
        70497 => X"1B",  -- 27
        70498 => X"17",  -- 23
        70499 => X"1C",  -- 28
        70500 => X"1F",  -- 31
        70501 => X"2C",  -- 44
        70502 => X"18",  -- 24
        70503 => X"19",  -- 25
        70504 => X"16",  -- 22
        70505 => X"1C",  -- 28
        70506 => X"19",  -- 25
        70507 => X"18",  -- 24
        70508 => X"1F",  -- 31
        70509 => X"1E",  -- 30
        70510 => X"15",  -- 21
        70511 => X"12",  -- 18
        70512 => X"17",  -- 23
        70513 => X"18",  -- 24
        70514 => X"1C",  -- 28
        70515 => X"23",  -- 35
        70516 => X"2A",  -- 42
        70517 => X"2D",  -- 45
        70518 => X"2B",  -- 43
        70519 => X"28",  -- 40
        70520 => X"30",  -- 48
        70521 => X"31",  -- 49
        70522 => X"33",  -- 51
        70523 => X"37",  -- 55
        70524 => X"35",  -- 53
        70525 => X"32",  -- 50
        70526 => X"36",  -- 54
        70527 => X"3E",  -- 62
        70528 => X"44",  -- 68
        70529 => X"3A",  -- 58
        70530 => X"2E",  -- 46
        70531 => X"2A",  -- 42
        70532 => X"2D",  -- 45
        70533 => X"33",  -- 51
        70534 => X"38",  -- 56
        70535 => X"3B",  -- 59
        70536 => X"44",  -- 68
        70537 => X"49",  -- 73
        70538 => X"35",  -- 53
        70539 => X"37",  -- 55
        70540 => X"40",  -- 64
        70541 => X"3A",  -- 58
        70542 => X"42",  -- 66
        70543 => X"48",  -- 72
        70544 => X"52",  -- 82
        70545 => X"3C",  -- 60
        70546 => X"42",  -- 66
        70547 => X"48",  -- 72
        70548 => X"61",  -- 97
        70549 => X"41",  -- 65
        70550 => X"4A",  -- 74
        70551 => X"3D",  -- 61
        70552 => X"3D",  -- 61
        70553 => X"3F",  -- 63
        70554 => X"3F",  -- 63
        70555 => X"3F",  -- 63
        70556 => X"3E",  -- 62
        70557 => X"3D",  -- 61
        70558 => X"3F",  -- 63
        70559 => X"40",  -- 64
        70560 => X"49",  -- 73
        70561 => X"3C",  -- 60
        70562 => X"4E",  -- 78
        70563 => X"48",  -- 72
        70564 => X"53",  -- 83
        70565 => X"57",  -- 87
        70566 => X"56",  -- 86
        70567 => X"5D",  -- 93
        70568 => X"4D",  -- 77
        70569 => X"41",  -- 65
        70570 => X"4A",  -- 74
        70571 => X"59",  -- 89
        70572 => X"5D",  -- 93
        70573 => X"52",  -- 82
        70574 => X"46",  -- 70
        70575 => X"4C",  -- 76
        70576 => X"55",  -- 85
        70577 => X"4C",  -- 76
        70578 => X"3A",  -- 58
        70579 => X"3F",  -- 63
        70580 => X"49",  -- 73
        70581 => X"49",  -- 73
        70582 => X"4F",  -- 79
        70583 => X"47",  -- 71
        70584 => X"67",  -- 103
        70585 => X"5B",  -- 91
        70586 => X"51",  -- 81
        70587 => X"47",  -- 71
        70588 => X"57",  -- 87
        70589 => X"63",  -- 99
        70590 => X"53",  -- 83
        70591 => X"50",  -- 80
        70592 => X"5B",  -- 91
        70593 => X"5E",  -- 94
        70594 => X"62",  -- 98
        70595 => X"60",  -- 96
        70596 => X"62",  -- 98
        70597 => X"69",  -- 105
        70598 => X"6E",  -- 110
        70599 => X"71",  -- 113
        70600 => X"6E",  -- 110
        70601 => X"72",  -- 114
        70602 => X"75",  -- 117
        70603 => X"6F",  -- 111
        70604 => X"64",  -- 100
        70605 => X"5A",  -- 90
        70606 => X"58",  -- 88
        70607 => X"58",  -- 88
        70608 => X"5B",  -- 91
        70609 => X"61",  -- 97
        70610 => X"62",  -- 98
        70611 => X"58",  -- 88
        70612 => X"54",  -- 84
        70613 => X"59",  -- 89
        70614 => X"5B",  -- 91
        70615 => X"58",  -- 88
        70616 => X"5C",  -- 92
        70617 => X"65",  -- 101
        70618 => X"70",  -- 112
        70619 => X"73",  -- 115
        70620 => X"6D",  -- 109
        70621 => X"6B",  -- 107
        70622 => X"71",  -- 113
        70623 => X"79",  -- 121
        70624 => X"91",  -- 145
        70625 => X"81",  -- 129
        70626 => X"6D",  -- 109
        70627 => X"7B",  -- 123
        70628 => X"87",  -- 135
        70629 => X"79",  -- 121
        70630 => X"76",  -- 118
        70631 => X"73",  -- 115
        70632 => X"66",  -- 102
        70633 => X"66",  -- 102
        70634 => X"68",  -- 104
        70635 => X"6C",  -- 108
        70636 => X"73",  -- 115
        70637 => X"78",  -- 120
        70638 => X"76",  -- 118
        70639 => X"70",  -- 112
        70640 => X"75",  -- 117
        70641 => X"75",  -- 117
        70642 => X"68",  -- 104
        70643 => X"6A",  -- 106
        70644 => X"73",  -- 115
        70645 => X"90",  -- 144
        70646 => X"83",  -- 131
        70647 => X"71",  -- 113
        70648 => X"72",  -- 114
        70649 => X"70",  -- 112
        70650 => X"69",  -- 105
        70651 => X"71",  -- 113
        70652 => X"8E",  -- 142
        70653 => X"7F",  -- 127
        70654 => X"7F",  -- 127
        70655 => X"78",  -- 120
        70656 => X"6B",  -- 107
        70657 => X"91",  -- 145
        70658 => X"8C",  -- 140
        70659 => X"68",  -- 104
        70660 => X"5D",  -- 93
        70661 => X"63",  -- 99
        70662 => X"76",  -- 118
        70663 => X"94",  -- 148
        70664 => X"8E",  -- 142
        70665 => X"87",  -- 135
        70666 => X"87",  -- 135
        70667 => X"8D",  -- 141
        70668 => X"97",  -- 151
        70669 => X"A2",  -- 162
        70670 => X"98",  -- 152
        70671 => X"8D",  -- 141
        70672 => X"91",  -- 145
        70673 => X"90",  -- 144
        70674 => X"9B",  -- 155
        70675 => X"7F",  -- 127
        70676 => X"80",  -- 128
        70677 => X"66",  -- 102
        70678 => X"7F",  -- 127
        70679 => X"99",  -- 153
        70680 => X"9F",  -- 159
        70681 => X"99",  -- 153
        70682 => X"9D",  -- 157
        70683 => X"A4",  -- 164
        70684 => X"A2",  -- 162
        70685 => X"95",  -- 149
        70686 => X"96",  -- 150
        70687 => X"A1",  -- 161
        70688 => X"94",  -- 148
        70689 => X"88",  -- 136
        70690 => X"8A",  -- 138
        70691 => X"82",  -- 130
        70692 => X"8E",  -- 142
        70693 => X"91",  -- 145
        70694 => X"74",  -- 116
        70695 => X"78",  -- 120
        70696 => X"95",  -- 149
        70697 => X"70",  -- 112
        70698 => X"6A",  -- 106
        70699 => X"67",  -- 103
        70700 => X"61",  -- 97
        70701 => X"53",  -- 83
        70702 => X"43",  -- 67
        70703 => X"4D",  -- 77
        70704 => X"63",  -- 99
        70705 => X"4B",  -- 75
        70706 => X"55",  -- 85
        70707 => X"55",  -- 85
        70708 => X"58",  -- 88
        70709 => X"3F",  -- 63
        70710 => X"3C",  -- 60
        70711 => X"35",  -- 53
        70712 => X"45",  -- 69
        70713 => X"58",  -- 88
        70714 => X"3E",  -- 62
        70715 => X"35",  -- 53
        70716 => X"4B",  -- 75
        70717 => X"65",  -- 101
        70718 => X"6F",  -- 111
        70719 => X"8F",  -- 143
        70720 => X"62",  -- 98
        70721 => X"60",  -- 96
        70722 => X"5E",  -- 94
        70723 => X"56",  -- 86
        70724 => X"52",  -- 82
        70725 => X"5F",  -- 95
        70726 => X"68",  -- 104
        70727 => X"62",  -- 98
        70728 => X"62",  -- 98
        70729 => X"64",  -- 100
        70730 => X"5A",  -- 90
        70731 => X"51",  -- 81
        70732 => X"54",  -- 84
        70733 => X"56",  -- 86
        70734 => X"50",  -- 80
        70735 => X"50",  -- 80
        70736 => X"4F",  -- 79
        70737 => X"52",  -- 82
        70738 => X"52",  -- 82
        70739 => X"51",  -- 81
        70740 => X"4D",  -- 77
        70741 => X"4E",  -- 78
        70742 => X"54",  -- 84
        70743 => X"59",  -- 89
        70744 => X"4E",  -- 78
        70745 => X"51",  -- 81
        70746 => X"57",  -- 87
        70747 => X"4E",  -- 78
        70748 => X"4F",  -- 79
        70749 => X"41",  -- 65
        70750 => X"68",  -- 104
        70751 => X"79",  -- 121
        70752 => X"4C",  -- 76
        70753 => X"45",  -- 69
        70754 => X"3B",  -- 59
        70755 => X"3B",  -- 59
        70756 => X"46",  -- 70
        70757 => X"4F",  -- 79
        70758 => X"4D",  -- 77
        70759 => X"46",  -- 70
        70760 => X"4D",  -- 77
        70761 => X"92",  -- 146
        70762 => X"7C",  -- 124
        70763 => X"3D",  -- 61
        70764 => X"43",  -- 67
        70765 => X"4A",  -- 74
        70766 => X"95",  -- 149
        70767 => X"43",  -- 67
        70768 => X"3E",  -- 62
        70769 => X"2A",  -- 42
        70770 => X"2E",  -- 46
        70771 => X"37",  -- 55
        70772 => X"3D",  -- 61
        70773 => X"22",  -- 34
        70774 => X"1E",  -- 30
        70775 => X"23",  -- 35
        70776 => X"1D",  -- 29
        70777 => X"18",  -- 24
        70778 => X"17",  -- 23
        70779 => X"2F",  -- 47
        70780 => X"3A",  -- 58
        70781 => X"2D",  -- 45
        70782 => X"28",  -- 40
        70783 => X"20",  -- 32
        70784 => X"25",  -- 37
        70785 => X"1E",  -- 30
        70786 => X"1C",  -- 28
        70787 => X"1B",  -- 27
        70788 => X"1D",  -- 29
        70789 => X"28",  -- 40
        70790 => X"2C",  -- 44
        70791 => X"20",  -- 32
        70792 => X"2A",  -- 42
        70793 => X"24",  -- 36
        70794 => X"32",  -- 50
        70795 => X"2E",  -- 46
        70796 => X"30",  -- 48
        70797 => X"1F",  -- 31
        70798 => X"25",  -- 37
        70799 => X"1E",  -- 30
        70800 => X"1D",  -- 29
        70801 => X"1A",  -- 26
        70802 => X"19",  -- 25
        70803 => X"1A",  -- 26
        70804 => X"1B",  -- 27
        70805 => X"1C",  -- 28
        70806 => X"21",  -- 33
        70807 => X"27",  -- 39
        70808 => X"2E",  -- 46
        70809 => X"25",  -- 37
        70810 => X"1E",  -- 30
        70811 => X"1F",  -- 31
        70812 => X"22",  -- 34
        70813 => X"1E",  -- 30
        70814 => X"16",  -- 22
        70815 => X"10",  -- 16
        70816 => X"10",  -- 16
        70817 => X"1F",  -- 31
        70818 => X"19",  -- 25
        70819 => X"1D",  -- 29
        70820 => X"1F",  -- 31
        70821 => X"2E",  -- 46
        70822 => X"1F",  -- 31
        70823 => X"1A",  -- 26
        70824 => X"16",  -- 22
        70825 => X"1A",  -- 26
        70826 => X"18",  -- 24
        70827 => X"18",  -- 24
        70828 => X"22",  -- 34
        70829 => X"23",  -- 35
        70830 => X"1A",  -- 26
        70831 => X"15",  -- 21
        70832 => X"1B",  -- 27
        70833 => X"1E",  -- 30
        70834 => X"23",  -- 35
        70835 => X"28",  -- 40
        70836 => X"2C",  -- 44
        70837 => X"30",  -- 48
        70838 => X"34",  -- 52
        70839 => X"38",  -- 56
        70840 => X"38",  -- 56
        70841 => X"36",  -- 54
        70842 => X"38",  -- 56
        70843 => X"3E",  -- 62
        70844 => X"3B",  -- 59
        70845 => X"35",  -- 53
        70846 => X"39",  -- 57
        70847 => X"45",  -- 69
        70848 => X"4B",  -- 75
        70849 => X"40",  -- 64
        70850 => X"36",  -- 54
        70851 => X"34",  -- 52
        70852 => X"38",  -- 56
        70853 => X"3C",  -- 60
        70854 => X"3F",  -- 63
        70855 => X"41",  -- 65
        70856 => X"49",  -- 73
        70857 => X"41",  -- 65
        70858 => X"2B",  -- 43
        70859 => X"3D",  -- 61
        70860 => X"3C",  -- 60
        70861 => X"2C",  -- 44
        70862 => X"3C",  -- 60
        70863 => X"3A",  -- 58
        70864 => X"64",  -- 100
        70865 => X"46",  -- 70
        70866 => X"38",  -- 56
        70867 => X"47",  -- 71
        70868 => X"63",  -- 99
        70869 => X"3C",  -- 60
        70870 => X"3C",  -- 60
        70871 => X"45",  -- 69
        70872 => X"42",  -- 66
        70873 => X"41",  -- 65
        70874 => X"40",  -- 64
        70875 => X"3F",  -- 63
        70876 => X"3F",  -- 63
        70877 => X"40",  -- 64
        70878 => X"41",  -- 65
        70879 => X"42",  -- 66
        70880 => X"4E",  -- 78
        70881 => X"3D",  -- 61
        70882 => X"3D",  -- 61
        70883 => X"3F",  -- 63
        70884 => X"54",  -- 84
        70885 => X"46",  -- 70
        70886 => X"53",  -- 83
        70887 => X"53",  -- 83
        70888 => X"6C",  -- 108
        70889 => X"56",  -- 86
        70890 => X"46",  -- 70
        70891 => X"46",  -- 70
        70892 => X"48",  -- 72
        70893 => X"44",  -- 68
        70894 => X"41",  -- 65
        70895 => X"44",  -- 68
        70896 => X"57",  -- 87
        70897 => X"5C",  -- 92
        70898 => X"53",  -- 83
        70899 => X"53",  -- 83
        70900 => X"56",  -- 86
        70901 => X"57",  -- 87
        70902 => X"5A",  -- 90
        70903 => X"4C",  -- 76
        70904 => X"64",  -- 100
        70905 => X"5D",  -- 93
        70906 => X"55",  -- 85
        70907 => X"4A",  -- 74
        70908 => X"58",  -- 88
        70909 => X"66",  -- 102
        70910 => X"5C",  -- 92
        70911 => X"5D",  -- 93
        70912 => X"59",  -- 89
        70913 => X"5E",  -- 94
        70914 => X"63",  -- 99
        70915 => X"63",  -- 99
        70916 => X"65",  -- 101
        70917 => X"69",  -- 105
        70918 => X"6D",  -- 109
        70919 => X"6E",  -- 110
        70920 => X"6F",  -- 111
        70921 => X"73",  -- 115
        70922 => X"74",  -- 116
        70923 => X"6F",  -- 111
        70924 => X"66",  -- 102
        70925 => X"5D",  -- 93
        70926 => X"5B",  -- 91
        70927 => X"5D",  -- 93
        70928 => X"61",  -- 97
        70929 => X"65",  -- 101
        70930 => X"64",  -- 100
        70931 => X"5F",  -- 95
        70932 => X"5C",  -- 92
        70933 => X"5B",  -- 91
        70934 => X"59",  -- 89
        70935 => X"58",  -- 88
        70936 => X"5D",  -- 93
        70937 => X"5C",  -- 92
        70938 => X"62",  -- 98
        70939 => X"70",  -- 112
        70940 => X"79",  -- 121
        70941 => X"7A",  -- 122
        70942 => X"7A",  -- 122
        70943 => X"7C",  -- 124
        70944 => X"89",  -- 137
        70945 => X"83",  -- 131
        70946 => X"74",  -- 116
        70947 => X"7A",  -- 122
        70948 => X"81",  -- 129
        70949 => X"7C",  -- 124
        70950 => X"7A",  -- 122
        70951 => X"6B",  -- 107
        70952 => X"67",  -- 103
        70953 => X"67",  -- 103
        70954 => X"63",  -- 99
        70955 => X"5E",  -- 94
        70956 => X"5A",  -- 90
        70957 => X"5C",  -- 92
        70958 => X"5F",  -- 95
        70959 => X"60",  -- 96
        70960 => X"6D",  -- 109
        70961 => X"6E",  -- 110
        70962 => X"63",  -- 99
        70963 => X"50",  -- 80
        70964 => X"70",  -- 112
        70965 => X"92",  -- 146
        70966 => X"98",  -- 152
        70967 => X"A9",  -- 169
        70968 => X"84",  -- 132
        70969 => X"70",  -- 112
        70970 => X"62",  -- 98
        70971 => X"65",  -- 101
        70972 => X"77",  -- 119
        70973 => X"6E",  -- 110
        70974 => X"74",  -- 116
        70975 => X"62",  -- 98
        70976 => X"5F",  -- 95
        70977 => X"7B",  -- 123
        70978 => X"90",  -- 144
        70979 => X"8F",  -- 143
        70980 => X"7B",  -- 123
        70981 => X"5C",  -- 92
        70982 => X"60",  -- 96
        70983 => X"83",  -- 131
        70984 => X"64",  -- 100
        70985 => X"5A",  -- 90
        70986 => X"84",  -- 132
        70987 => X"74",  -- 116
        70988 => X"98",  -- 152
        70989 => X"8A",  -- 138
        70990 => X"95",  -- 149
        70991 => X"7E",  -- 126
        70992 => X"8E",  -- 142
        70993 => X"8D",  -- 141
        70994 => X"6F",  -- 111
        70995 => X"7B",  -- 123
        70996 => X"82",  -- 130
        70997 => X"78",  -- 120
        70998 => X"96",  -- 150
        70999 => X"A5",  -- 165
        71000 => X"99",  -- 153
        71001 => X"92",  -- 146
        71002 => X"92",  -- 146
        71003 => X"91",  -- 145
        71004 => X"9A",  -- 154
        71005 => X"94",  -- 148
        71006 => X"93",  -- 147
        71007 => X"8F",  -- 143
        71008 => X"7C",  -- 124
        71009 => X"81",  -- 129
        71010 => X"8A",  -- 138
        71011 => X"8F",  -- 143
        71012 => X"8F",  -- 143
        71013 => X"7A",  -- 122
        71014 => X"6A",  -- 106
        71015 => X"83",  -- 131
        71016 => X"8F",  -- 143
        71017 => X"65",  -- 101
        71018 => X"60",  -- 96
        71019 => X"5D",  -- 93
        71020 => X"6D",  -- 109
        71021 => X"5B",  -- 91
        71022 => X"4C",  -- 76
        71023 => X"6A",  -- 106
        71024 => X"5F",  -- 95
        71025 => X"63",  -- 99
        71026 => X"6B",  -- 107
        71027 => X"6F",  -- 111
        71028 => X"52",  -- 82
        71029 => X"54",  -- 84
        71030 => X"42",  -- 66
        71031 => X"44",  -- 68
        71032 => X"3E",  -- 62
        71033 => X"3E",  -- 62
        71034 => X"3B",  -- 59
        71035 => X"35",  -- 53
        71036 => X"33",  -- 51
        71037 => X"5B",  -- 91
        71038 => X"83",  -- 131
        71039 => X"8C",  -- 140
        71040 => X"5A",  -- 90
        71041 => X"57",  -- 87
        71042 => X"59",  -- 89
        71043 => X"59",  -- 89
        71044 => X"4F",  -- 79
        71045 => X"51",  -- 81
        71046 => X"5B",  -- 91
        71047 => X"5E",  -- 94
        71048 => X"54",  -- 84
        71049 => X"5A",  -- 90
        71050 => X"59",  -- 89
        71051 => X"5B",  -- 91
        71052 => X"64",  -- 100
        71053 => X"5F",  -- 95
        71054 => X"52",  -- 82
        71055 => X"4A",  -- 74
        71056 => X"4C",  -- 76
        71057 => X"51",  -- 81
        71058 => X"59",  -- 89
        71059 => X"5A",  -- 90
        71060 => X"57",  -- 87
        71061 => X"56",  -- 86
        71062 => X"5A",  -- 90
        71063 => X"5D",  -- 93
        71064 => X"4B",  -- 75
        71065 => X"4E",  -- 78
        71066 => X"50",  -- 80
        71067 => X"51",  -- 81
        71068 => X"4C",  -- 76
        71069 => X"55",  -- 85
        71070 => X"72",  -- 114
        71071 => X"6E",  -- 110
        71072 => X"5B",  -- 91
        71073 => X"45",  -- 69
        71074 => X"37",  -- 55
        71075 => X"3A",  -- 58
        71076 => X"43",  -- 67
        71077 => X"44",  -- 68
        71078 => X"42",  -- 66
        71079 => X"45",  -- 69
        71080 => X"56",  -- 86
        71081 => X"87",  -- 135
        71082 => X"7E",  -- 126
        71083 => X"51",  -- 81
        71084 => X"44",  -- 68
        71085 => X"58",  -- 88
        71086 => X"83",  -- 131
        71087 => X"39",  -- 57
        71088 => X"46",  -- 70
        71089 => X"38",  -- 56
        71090 => X"39",  -- 57
        71091 => X"38",  -- 56
        71092 => X"3D",  -- 61
        71093 => X"2B",  -- 43
        71094 => X"29",  -- 41
        71095 => X"29",  -- 41
        71096 => X"2C",  -- 44
        71097 => X"24",  -- 36
        71098 => X"17",  -- 23
        71099 => X"2A",  -- 42
        71100 => X"2E",  -- 46
        71101 => X"1E",  -- 30
        71102 => X"20",  -- 32
        71103 => X"1A",  -- 26
        71104 => X"21",  -- 33
        71105 => X"1E",  -- 30
        71106 => X"22",  -- 34
        71107 => X"26",  -- 38
        71108 => X"24",  -- 36
        71109 => X"28",  -- 40
        71110 => X"28",  -- 40
        71111 => X"21",  -- 33
        71112 => X"23",  -- 35
        71113 => X"23",  -- 35
        71114 => X"2C",  -- 44
        71115 => X"2A",  -- 42
        71116 => X"2A",  -- 42
        71117 => X"1E",  -- 30
        71118 => X"20",  -- 32
        71119 => X"1F",  -- 31
        71120 => X"1F",  -- 31
        71121 => X"1A",  -- 26
        71122 => X"17",  -- 23
        71123 => X"1A",  -- 26
        71124 => X"1C",  -- 28
        71125 => X"1D",  -- 29
        71126 => X"1E",  -- 30
        71127 => X"21",  -- 33
        71128 => X"2C",  -- 44
        71129 => X"26",  -- 38
        71130 => X"22",  -- 34
        71131 => X"23",  -- 35
        71132 => X"23",  -- 35
        71133 => X"1F",  -- 31
        71134 => X"1C",  -- 28
        71135 => X"1C",  -- 28
        71136 => X"16",  -- 22
        71137 => X"24",  -- 36
        71138 => X"19",  -- 25
        71139 => X"1E",  -- 30
        71140 => X"1D",  -- 29
        71141 => X"25",  -- 37
        71142 => X"1A",  -- 26
        71143 => X"16",  -- 22
        71144 => X"16",  -- 22
        71145 => X"1B",  -- 27
        71146 => X"19",  -- 25
        71147 => X"1B",  -- 27
        71148 => X"29",  -- 41
        71149 => X"2C",  -- 44
        71150 => X"22",  -- 34
        71151 => X"1C",  -- 28
        71152 => X"23",  -- 35
        71153 => X"25",  -- 37
        71154 => X"27",  -- 39
        71155 => X"28",  -- 40
        71156 => X"2C",  -- 44
        71157 => X"33",  -- 51
        71158 => X"3B",  -- 59
        71159 => X"41",  -- 65
        71160 => X"3D",  -- 61
        71161 => X"35",  -- 53
        71162 => X"35",  -- 53
        71163 => X"3C",  -- 60
        71164 => X"3A",  -- 58
        71165 => X"32",  -- 50
        71166 => X"35",  -- 53
        71167 => X"3F",  -- 63
        71168 => X"40",  -- 64
        71169 => X"3B",  -- 59
        71170 => X"37",  -- 55
        71171 => X"38",  -- 56
        71172 => X"3A",  -- 58
        71173 => X"3B",  -- 59
        71174 => X"3F",  -- 63
        71175 => X"45",  -- 69
        71176 => X"4B",  -- 75
        71177 => X"3C",  -- 60
        71178 => X"3D",  -- 61
        71179 => X"43",  -- 67
        71180 => X"34",  -- 52
        71181 => X"31",  -- 49
        71182 => X"3A",  -- 58
        71183 => X"31",  -- 49
        71184 => X"61",  -- 97
        71185 => X"52",  -- 82
        71186 => X"37",  -- 55
        71187 => X"44",  -- 68
        71188 => X"5D",  -- 93
        71189 => X"3C",  -- 60
        71190 => X"32",  -- 50
        71191 => X"45",  -- 69
        71192 => X"42",  -- 66
        71193 => X"3F",  -- 63
        71194 => X"3F",  -- 63
        71195 => X"41",  -- 65
        71196 => X"46",  -- 70
        71197 => X"4A",  -- 74
        71198 => X"4C",  -- 76
        71199 => X"4D",  -- 77
        71200 => X"4E",  -- 78
        71201 => X"46",  -- 70
        71202 => X"3E",  -- 62
        71203 => X"40",  -- 64
        71204 => X"46",  -- 70
        71205 => X"3C",  -- 60
        71206 => X"42",  -- 66
        71207 => X"52",  -- 82
        71208 => X"61",  -- 97
        71209 => X"59",  -- 89
        71210 => X"4F",  -- 79
        71211 => X"52",  -- 82
        71212 => X"54",  -- 84
        71213 => X"4E",  -- 78
        71214 => X"48",  -- 72
        71215 => X"41",  -- 65
        71216 => X"52",  -- 82
        71217 => X"5B",  -- 91
        71218 => X"58",  -- 88
        71219 => X"5C",  -- 92
        71220 => X"5C",  -- 92
        71221 => X"55",  -- 85
        71222 => X"55",  -- 85
        71223 => X"47",  -- 71
        71224 => X"4E",  -- 78
        71225 => X"50",  -- 80
        71226 => X"50",  -- 80
        71227 => X"47",  -- 71
        71228 => X"51",  -- 81
        71229 => X"5F",  -- 95
        71230 => X"57",  -- 87
        71231 => X"5B",  -- 91
        71232 => X"58",  -- 88
        71233 => X"5D",  -- 93
        71234 => X"62",  -- 98
        71235 => X"63",  -- 99
        71236 => X"65",  -- 101
        71237 => X"69",  -- 105
        71238 => X"6C",  -- 108
        71239 => X"6B",  -- 107
        71240 => X"6B",  -- 107
        71241 => X"6E",  -- 110
        71242 => X"70",  -- 112
        71243 => X"6D",  -- 109
        71244 => X"66",  -- 102
        71245 => X"62",  -- 98
        71246 => X"5F",  -- 95
        71247 => X"60",  -- 96
        71248 => X"61",  -- 97
        71249 => X"5E",  -- 94
        71250 => X"5D",  -- 93
        71251 => X"62",  -- 98
        71252 => X"64",  -- 100
        71253 => X"60",  -- 96
        71254 => X"5C",  -- 92
        71255 => X"59",  -- 89
        71256 => X"60",  -- 96
        71257 => X"62",  -- 98
        71258 => X"68",  -- 104
        71259 => X"70",  -- 112
        71260 => X"7B",  -- 123
        71261 => X"80",  -- 128
        71262 => X"7C",  -- 124
        71263 => X"76",  -- 118
        71264 => X"74",  -- 116
        71265 => X"7A",  -- 122
        71266 => X"76",  -- 118
        71267 => X"7A",  -- 122
        71268 => X"7B",  -- 123
        71269 => X"7A",  -- 122
        71270 => X"79",  -- 121
        71271 => X"65",  -- 101
        71272 => X"66",  -- 102
        71273 => X"61",  -- 97
        71274 => X"5A",  -- 90
        71275 => X"56",  -- 86
        71276 => X"5F",  -- 95
        71277 => X"69",  -- 105
        71278 => X"6B",  -- 107
        71279 => X"66",  -- 102
        71280 => X"59",  -- 89
        71281 => X"73",  -- 115
        71282 => X"6C",  -- 108
        71283 => X"5B",  -- 91
        71284 => X"8A",  -- 138
        71285 => X"81",  -- 129
        71286 => X"83",  -- 131
        71287 => X"8F",  -- 143
        71288 => X"81",  -- 129
        71289 => X"72",  -- 114
        71290 => X"74",  -- 116
        71291 => X"76",  -- 118
        71292 => X"74",  -- 116
        71293 => X"6C",  -- 108
        71294 => X"7E",  -- 126
        71295 => X"69",  -- 105
        71296 => X"7A",  -- 122
        71297 => X"69",  -- 105
        71298 => X"6A",  -- 106
        71299 => X"7D",  -- 125
        71300 => X"76",  -- 118
        71301 => X"5D",  -- 93
        71302 => X"63",  -- 99
        71303 => X"84",  -- 132
        71304 => X"5D",  -- 93
        71305 => X"4E",  -- 78
        71306 => X"7F",  -- 127
        71307 => X"7C",  -- 124
        71308 => X"91",  -- 145
        71309 => X"7F",  -- 127
        71310 => X"86",  -- 134
        71311 => X"7D",  -- 125
        71312 => X"83",  -- 131
        71313 => X"87",  -- 135
        71314 => X"65",  -- 101
        71315 => X"85",  -- 133
        71316 => X"95",  -- 149
        71317 => X"96",  -- 150
        71318 => X"99",  -- 153
        71319 => X"8F",  -- 143
        71320 => X"89",  -- 137
        71321 => X"9B",  -- 155
        71322 => X"A9",  -- 169
        71323 => X"8E",  -- 142
        71324 => X"86",  -- 134
        71325 => X"7B",  -- 123
        71326 => X"80",  -- 128
        71327 => X"76",  -- 118
        71328 => X"7C",  -- 124
        71329 => X"6D",  -- 109
        71330 => X"5C",  -- 92
        71331 => X"7B",  -- 123
        71332 => X"94",  -- 148
        71333 => X"79",  -- 121
        71334 => X"6A",  -- 106
        71335 => X"7E",  -- 126
        71336 => X"74",  -- 116
        71337 => X"61",  -- 97
        71338 => X"5E",  -- 94
        71339 => X"47",  -- 71
        71340 => X"69",  -- 105
        71341 => X"67",  -- 103
        71342 => X"51",  -- 81
        71343 => X"69",  -- 105
        71344 => X"7B",  -- 123
        71345 => X"76",  -- 118
        71346 => X"73",  -- 115
        71347 => X"66",  -- 102
        71348 => X"48",  -- 72
        71349 => X"5A",  -- 90
        71350 => X"55",  -- 85
        71351 => X"60",  -- 96
        71352 => X"46",  -- 70
        71353 => X"2F",  -- 47
        71354 => X"32",  -- 50
        71355 => X"3F",  -- 63
        71356 => X"3B",  -- 59
        71357 => X"43",  -- 67
        71358 => X"6D",  -- 109
        71359 => X"91",  -- 145
        71360 => X"65",  -- 101
        71361 => X"60",  -- 96
        71362 => X"68",  -- 104
        71363 => X"6C",  -- 108
        71364 => X"5D",  -- 93
        71365 => X"51",  -- 81
        71366 => X"58",  -- 88
        71367 => X"5F",  -- 95
        71368 => X"60",  -- 96
        71369 => X"63",  -- 99
        71370 => X"5F",  -- 95
        71371 => X"5E",  -- 94
        71372 => X"65",  -- 101
        71373 => X"5F",  -- 95
        71374 => X"51",  -- 81
        71375 => X"4D",  -- 77
        71376 => X"4C",  -- 76
        71377 => X"53",  -- 83
        71378 => X"59",  -- 89
        71379 => X"5B",  -- 91
        71380 => X"58",  -- 88
        71381 => X"57",  -- 87
        71382 => X"5A",  -- 90
        71383 => X"5D",  -- 93
        71384 => X"46",  -- 70
        71385 => X"40",  -- 64
        71386 => X"32",  -- 50
        71387 => X"42",  -- 66
        71388 => X"3E",  -- 62
        71389 => X"64",  -- 100
        71390 => X"73",  -- 115
        71391 => X"59",  -- 89
        71392 => X"61",  -- 97
        71393 => X"4D",  -- 77
        71394 => X"3C",  -- 60
        71395 => X"3B",  -- 59
        71396 => X"44",  -- 68
        71397 => X"46",  -- 70
        71398 => X"40",  -- 64
        71399 => X"3D",  -- 61
        71400 => X"59",  -- 89
        71401 => X"6D",  -- 109
        71402 => X"61",  -- 97
        71403 => X"5B",  -- 91
        71404 => X"2F",  -- 47
        71405 => X"61",  -- 97
        71406 => X"6A",  -- 106
        71407 => X"4A",  -- 74
        71408 => X"44",  -- 68
        71409 => X"43",  -- 67
        71410 => X"3F",  -- 63
        71411 => X"3C",  -- 60
        71412 => X"38",  -- 56
        71413 => X"32",  -- 50
        71414 => X"2A",  -- 42
        71415 => X"24",  -- 36
        71416 => X"27",  -- 39
        71417 => X"2B",  -- 43
        71418 => X"23",  -- 35
        71419 => X"2E",  -- 46
        71420 => X"2B",  -- 43
        71421 => X"18",  -- 24
        71422 => X"24",  -- 36
        71423 => X"26",  -- 38
        71424 => X"25",  -- 37
        71425 => X"22",  -- 34
        71426 => X"2A",  -- 42
        71427 => X"2E",  -- 46
        71428 => X"25",  -- 37
        71429 => X"1E",  -- 30
        71430 => X"1C",  -- 28
        71431 => X"16",  -- 22
        71432 => X"16",  -- 22
        71433 => X"19",  -- 25
        71434 => X"21",  -- 33
        71435 => X"23",  -- 35
        71436 => X"21",  -- 33
        71437 => X"1C",  -- 28
        71438 => X"1D",  -- 29
        71439 => X"20",  -- 32
        71440 => X"1F",  -- 31
        71441 => X"1A",  -- 26
        71442 => X"1A",  -- 26
        71443 => X"21",  -- 33
        71444 => X"27",  -- 39
        71445 => X"23",  -- 35
        71446 => X"1C",  -- 28
        71447 => X"18",  -- 24
        71448 => X"1C",  -- 28
        71449 => X"1C",  -- 28
        71450 => X"20",  -- 32
        71451 => X"25",  -- 37
        71452 => X"24",  -- 36
        71453 => X"1F",  -- 31
        71454 => X"1E",  -- 30
        71455 => X"23",  -- 35
        71456 => X"19",  -- 25
        71457 => X"23",  -- 35
        71458 => X"14",  -- 20
        71459 => X"1B",  -- 27
        71460 => X"15",  -- 21
        71461 => X"13",  -- 19
        71462 => X"09",  -- 9
        71463 => X"09",  -- 9
        71464 => X"13",  -- 19
        71465 => X"18",  -- 24
        71466 => X"17",  -- 23
        71467 => X"1B",  -- 27
        71468 => X"2A",  -- 42
        71469 => X"2C",  -- 44
        71470 => X"23",  -- 35
        71471 => X"1B",  -- 27
        71472 => X"2C",  -- 44
        71473 => X"2C",  -- 44
        71474 => X"2B",  -- 43
        71475 => X"2A",  -- 42
        71476 => X"2C",  -- 44
        71477 => X"30",  -- 48
        71478 => X"36",  -- 54
        71479 => X"3B",  -- 59
        71480 => X"40",  -- 64
        71481 => X"32",  -- 50
        71482 => X"2D",  -- 45
        71483 => X"34",  -- 52
        71484 => X"34",  -- 52
        71485 => X"2B",  -- 43
        71486 => X"29",  -- 41
        71487 => X"30",  -- 48
        71488 => X"32",  -- 50
        71489 => X"32",  -- 50
        71490 => X"35",  -- 53
        71491 => X"38",  -- 56
        71492 => X"36",  -- 54
        71493 => X"35",  -- 53
        71494 => X"3D",  -- 61
        71495 => X"47",  -- 71
        71496 => X"45",  -- 69
        71497 => X"3D",  -- 61
        71498 => X"5A",  -- 90
        71499 => X"48",  -- 72
        71500 => X"30",  -- 48
        71501 => X"4A",  -- 74
        71502 => X"4B",  -- 75
        71503 => X"37",  -- 55
        71504 => X"41",  -- 65
        71505 => X"53",  -- 83
        71506 => X"36",  -- 54
        71507 => X"3B",  -- 59
        71508 => X"57",  -- 87
        71509 => X"4A",  -- 74
        71510 => X"39",  -- 57
        71511 => X"45",  -- 69
        71512 => X"47",  -- 71
        71513 => X"44",  -- 68
        71514 => X"40",  -- 64
        71515 => X"41",  -- 65
        71516 => X"47",  -- 71
        71517 => X"4D",  -- 77
        71518 => X"4F",  -- 79
        71519 => X"50",  -- 80
        71520 => X"47",  -- 71
        71521 => X"4F",  -- 79
        71522 => X"4C",  -- 76
        71523 => X"4C",  -- 76
        71524 => X"3F",  -- 63
        71525 => X"42",  -- 66
        71526 => X"40",  -- 64
        71527 => X"6B",  -- 107
        71528 => X"49",  -- 73
        71529 => X"51",  -- 81
        71530 => X"54",  -- 84
        71531 => X"5D",  -- 93
        71532 => X"60",  -- 96
        71533 => X"5D",  -- 93
        71534 => X"5F",  -- 95
        71535 => X"5C",  -- 92
        71536 => X"5E",  -- 94
        71537 => X"59",  -- 89
        71538 => X"4C",  -- 76
        71539 => X"54",  -- 84
        71540 => X"5A",  -- 90
        71541 => X"57",  -- 87
        71542 => X"5A",  -- 90
        71543 => X"53",  -- 83
        71544 => X"4F",  -- 79
        71545 => X"59",  -- 89
        71546 => X"61",  -- 97
        71547 => X"58",  -- 88
        71548 => X"5E",  -- 94
        71549 => X"66",  -- 102
        71550 => X"5A",  -- 90
        71551 => X"5B",  -- 91
        71552 => X"5E",  -- 94
        71553 => X"62",  -- 98
        71554 => X"67",  -- 103
        71555 => X"67",  -- 103
        71556 => X"69",  -- 105
        71557 => X"6F",  -- 111
        71558 => X"70",  -- 112
        71559 => X"6F",  -- 111
        71560 => X"68",  -- 104
        71561 => X"69",  -- 105
        71562 => X"6C",  -- 108
        71563 => X"6A",  -- 106
        71564 => X"67",  -- 103
        71565 => X"64",  -- 100
        71566 => X"63",  -- 99
        71567 => X"63",  -- 99
        71568 => X"5E",  -- 94
        71569 => X"53",  -- 83
        71570 => X"51",  -- 81
        71571 => X"5F",  -- 95
        71572 => X"68",  -- 104
        71573 => X"65",  -- 101
        71574 => X"5C",  -- 92
        71575 => X"57",  -- 87
        71576 => X"62",  -- 98
        71577 => X"70",  -- 112
        71578 => X"78",  -- 120
        71579 => X"75",  -- 117
        71580 => X"73",  -- 115
        71581 => X"79",  -- 121
        71582 => X"78",  -- 120
        71583 => X"6E",  -- 110
        71584 => X"6D",  -- 109
        71585 => X"71",  -- 113
        71586 => X"73",  -- 115
        71587 => X"7F",  -- 127
        71588 => X"78",  -- 120
        71589 => X"6D",  -- 109
        71590 => X"6B",  -- 107
        71591 => X"5B",  -- 91
        71592 => X"54",  -- 84
        71593 => X"56",  -- 86
        71594 => X"57",  -- 87
        71595 => X"58",  -- 88
        71596 => X"62",  -- 98
        71597 => X"6D",  -- 109
        71598 => X"71",  -- 113
        71599 => X"6E",  -- 110
        71600 => X"6A",  -- 106
        71601 => X"8F",  -- 143
        71602 => X"72",  -- 114
        71603 => X"5E",  -- 94
        71604 => X"94",  -- 148
        71605 => X"67",  -- 103
        71606 => X"69",  -- 105
        71607 => X"66",  -- 102
        71608 => X"61",  -- 97
        71609 => X"66",  -- 102
        71610 => X"85",  -- 133
        71611 => X"8B",  -- 139
        71612 => X"76",  -- 118
        71613 => X"68",  -- 104
        71614 => X"84",  -- 132
        71615 => X"71",  -- 113
        71616 => X"6E",  -- 110
        71617 => X"6D",  -- 109
        71618 => X"6D",  -- 109
        71619 => X"69",  -- 105
        71620 => X"6C",  -- 108
        71621 => X"7D",  -- 125
        71622 => X"86",  -- 134
        71623 => X"7E",  -- 126
        71624 => X"7E",  -- 126
        71625 => X"64",  -- 100
        71626 => X"71",  -- 113
        71627 => X"87",  -- 135
        71628 => X"74",  -- 116
        71629 => X"7A",  -- 122
        71630 => X"70",  -- 112
        71631 => X"81",  -- 129
        71632 => X"7A",  -- 122
        71633 => X"91",  -- 145
        71634 => X"8E",  -- 142
        71635 => X"97",  -- 151
        71636 => X"9F",  -- 159
        71637 => X"96",  -- 150
        71638 => X"98",  -- 152
        71639 => X"8D",  -- 141
        71640 => X"97",  -- 151
        71641 => X"8D",  -- 141
        71642 => X"99",  -- 153
        71643 => X"9C",  -- 156
        71644 => X"A8",  -- 168
        71645 => X"8D",  -- 141
        71646 => X"7E",  -- 126
        71647 => X"6E",  -- 110
        71648 => X"6E",  -- 110
        71649 => X"5B",  -- 91
        71650 => X"3D",  -- 61
        71651 => X"60",  -- 96
        71652 => X"75",  -- 117
        71653 => X"4F",  -- 79
        71654 => X"52",  -- 82
        71655 => X"74",  -- 116
        71656 => X"87",  -- 135
        71657 => X"6F",  -- 111
        71658 => X"67",  -- 103
        71659 => X"52",  -- 82
        71660 => X"79",  -- 121
        71661 => X"66",  -- 102
        71662 => X"47",  -- 71
        71663 => X"68",  -- 104
        71664 => X"6A",  -- 106
        71665 => X"63",  -- 99
        71666 => X"81",  -- 129
        71667 => X"74",  -- 116
        71668 => X"77",  -- 119
        71669 => X"6F",  -- 111
        71670 => X"60",  -- 96
        71671 => X"53",  -- 83
        71672 => X"63",  -- 99
        71673 => X"59",  -- 89
        71674 => X"45",  -- 69
        71675 => X"42",  -- 66
        71676 => X"4A",  -- 74
        71677 => X"31",  -- 49
        71678 => X"40",  -- 64
        71679 => X"7F",  -- 127
        71680 => X"5C",  -- 92
        71681 => X"5A",  -- 90
        71682 => X"62",  -- 98
        71683 => X"6C",  -- 108
        71684 => X"66",  -- 102
        71685 => X"59",  -- 89
        71686 => X"5B",  -- 91
        71687 => X"6A",  -- 106
        71688 => X"62",  -- 98
        71689 => X"54",  -- 84
        71690 => X"52",  -- 82
        71691 => X"5D",  -- 93
        71692 => X"61",  -- 97
        71693 => X"55",  -- 85
        71694 => X"4A",  -- 74
        71695 => X"49",  -- 73
        71696 => X"44",  -- 68
        71697 => X"49",  -- 73
        71698 => X"53",  -- 83
        71699 => X"5E",  -- 94
        71700 => X"64",  -- 100
        71701 => X"62",  -- 98
        71702 => X"5C",  -- 92
        71703 => X"58",  -- 88
        71704 => X"54",  -- 84
        71705 => X"4A",  -- 74
        71706 => X"38",  -- 56
        71707 => X"41",  -- 65
        71708 => X"44",  -- 68
        71709 => X"7A",  -- 122
        71710 => X"44",  -- 68
        71711 => X"5A",  -- 90
        71712 => X"5B",  -- 91
        71713 => X"40",  -- 64
        71714 => X"3F",  -- 63
        71715 => X"3E",  -- 62
        71716 => X"3F",  -- 63
        71717 => X"45",  -- 69
        71718 => X"40",  -- 64
        71719 => X"44",  -- 68
        71720 => X"5E",  -- 94
        71721 => X"50",  -- 80
        71722 => X"31",  -- 49
        71723 => X"44",  -- 68
        71724 => X"45",  -- 69
        71725 => X"5A",  -- 90
        71726 => X"63",  -- 99
        71727 => X"49",  -- 73
        71728 => X"41",  -- 65
        71729 => X"36",  -- 54
        71730 => X"27",  -- 39
        71731 => X"34",  -- 52
        71732 => X"29",  -- 41
        71733 => X"2B",  -- 43
        71734 => X"1E",  -- 30
        71735 => X"25",  -- 37
        71736 => X"1E",  -- 30
        71737 => X"20",  -- 32
        71738 => X"24",  -- 36
        71739 => X"25",  -- 37
        71740 => X"1F",  -- 31
        71741 => X"18",  -- 24
        71742 => X"18",  -- 24
        71743 => X"1D",  -- 29
        71744 => X"1D",  -- 29
        71745 => X"27",  -- 39
        71746 => X"2D",  -- 45
        71747 => X"2A",  -- 42
        71748 => X"27",  -- 39
        71749 => X"25",  -- 37
        71750 => X"1D",  -- 29
        71751 => X"13",  -- 19
        71752 => X"13",  -- 19
        71753 => X"1B",  -- 27
        71754 => X"23",  -- 35
        71755 => X"24",  -- 36
        71756 => X"1E",  -- 30
        71757 => X"1B",  -- 27
        71758 => X"1F",  -- 31
        71759 => X"25",  -- 37
        71760 => X"1F",  -- 31
        71761 => X"14",  -- 20
        71762 => X"16",  -- 22
        71763 => X"21",  -- 33
        71764 => X"23",  -- 35
        71765 => X"20",  -- 32
        71766 => X"19",  -- 25
        71767 => X"0D",  -- 13
        71768 => X"10",  -- 16
        71769 => X"18",  -- 24
        71770 => X"1F",  -- 31
        71771 => X"20",  -- 32
        71772 => X"20",  -- 32
        71773 => X"20",  -- 32
        71774 => X"1F",  -- 31
        71775 => X"1C",  -- 28
        71776 => X"1A",  -- 26
        71777 => X"19",  -- 25
        71778 => X"1A",  -- 26
        71779 => X"18",  -- 24
        71780 => X"12",  -- 18
        71781 => X"0C",  -- 12
        71782 => X"0E",  -- 14
        71783 => X"14",  -- 20
        71784 => X"1E",  -- 30
        71785 => X"16",  -- 22
        71786 => X"15",  -- 21
        71787 => X"1D",  -- 29
        71788 => X"22",  -- 34
        71789 => X"1E",  -- 30
        71790 => X"18",  -- 24
        71791 => X"17",  -- 23
        71792 => X"25",  -- 37
        71793 => X"24",  -- 36
        71794 => X"2C",  -- 44
        71795 => X"2E",  -- 46
        71796 => X"27",  -- 39
        71797 => X"28",  -- 40
        71798 => X"34",  -- 52
        71799 => X"39",  -- 57
        71800 => X"34",  -- 52
        71801 => X"2D",  -- 45
        71802 => X"28",  -- 40
        71803 => X"2A",  -- 42
        71804 => X"2C",  -- 44
        71805 => X"2A",  -- 42
        71806 => X"2A",  -- 42
        71807 => X"2D",  -- 45
        71808 => X"3C",  -- 60
        71809 => X"31",  -- 49
        71810 => X"29",  -- 41
        71811 => X"2C",  -- 44
        71812 => X"32",  -- 50
        71813 => X"38",  -- 56
        71814 => X"3F",  -- 63
        71815 => X"47",  -- 71
        71816 => X"50",  -- 80
        71817 => X"49",  -- 73
        71818 => X"3E",  -- 62
        71819 => X"38",  -- 56
        71820 => X"35",  -- 53
        71821 => X"38",  -- 56
        71822 => X"3A",  -- 58
        71823 => X"3C",  -- 60
        71824 => X"3A",  -- 58
        71825 => X"57",  -- 87
        71826 => X"34",  -- 52
        71827 => X"40",  -- 64
        71828 => X"55",  -- 85
        71829 => X"46",  -- 70
        71830 => X"4C",  -- 76
        71831 => X"3C",  -- 60
        71832 => X"3E",  -- 62
        71833 => X"3B",  -- 59
        71834 => X"46",  -- 70
        71835 => X"47",  -- 71
        71836 => X"3B",  -- 59
        71837 => X"49",  -- 73
        71838 => X"52",  -- 82
        71839 => X"3A",  -- 58
        71840 => X"4A",  -- 74
        71841 => X"47",  -- 71
        71842 => X"41",  -- 65
        71843 => X"50",  -- 80
        71844 => X"58",  -- 88
        71845 => X"54",  -- 84
        71846 => X"5B",  -- 91
        71847 => X"58",  -- 88
        71848 => X"4C",  -- 76
        71849 => X"5A",  -- 90
        71850 => X"64",  -- 100
        71851 => X"66",  -- 102
        71852 => X"66",  -- 102
        71853 => X"6A",  -- 106
        71854 => X"71",  -- 113
        71855 => X"73",  -- 115
        71856 => X"72",  -- 114
        71857 => X"68",  -- 104
        71858 => X"61",  -- 97
        71859 => X"61",  -- 97
        71860 => X"62",  -- 98
        71861 => X"5C",  -- 92
        71862 => X"50",  -- 80
        71863 => X"49",  -- 73
        71864 => X"5C",  -- 92
        71865 => X"5D",  -- 93
        71866 => X"5C",  -- 92
        71867 => X"61",  -- 97
        71868 => X"62",  -- 98
        71869 => X"58",  -- 88
        71870 => X"56",  -- 86
        71871 => X"60",  -- 96
        71872 => X"61",  -- 97
        71873 => X"67",  -- 103
        71874 => X"59",  -- 89
        71875 => X"50",  -- 80
        71876 => X"60",  -- 96
        71877 => X"66",  -- 102
        71878 => X"64",  -- 100
        71879 => X"6C",  -- 108
        71880 => X"63",  -- 99
        71881 => X"6B",  -- 107
        71882 => X"6A",  -- 106
        71883 => X"64",  -- 100
        71884 => X"67",  -- 103
        71885 => X"65",  -- 101
        71886 => X"60",  -- 96
        71887 => X"62",  -- 98
        71888 => X"59",  -- 89
        71889 => X"5B",  -- 91
        71890 => X"5C",  -- 92
        71891 => X"5C",  -- 92
        71892 => X"5E",  -- 94
        71893 => X"62",  -- 98
        71894 => X"66",  -- 102
        71895 => X"66",  -- 102
        71896 => X"74",  -- 116
        71897 => X"70",  -- 112
        71898 => X"63",  -- 99
        71899 => X"66",  -- 102
        71900 => X"6D",  -- 109
        71901 => X"74",  -- 116
        71902 => X"5C",  -- 92
        71903 => X"68",  -- 104
        71904 => X"7B",  -- 123
        71905 => X"71",  -- 113
        71906 => X"70",  -- 112
        71907 => X"78",  -- 120
        71908 => X"76",  -- 118
        71909 => X"67",  -- 103
        71910 => X"5D",  -- 93
        71911 => X"5F",  -- 95
        71912 => X"53",  -- 83
        71913 => X"4C",  -- 76
        71914 => X"49",  -- 73
        71915 => X"4E",  -- 78
        71916 => X"5D",  -- 93
        71917 => X"6B",  -- 107
        71918 => X"71",  -- 113
        71919 => X"71",  -- 113
        71920 => X"7F",  -- 127
        71921 => X"73",  -- 115
        71922 => X"7C",  -- 124
        71923 => X"8D",  -- 141
        71924 => X"8A",  -- 138
        71925 => X"7D",  -- 125
        71926 => X"63",  -- 99
        71927 => X"42",  -- 66
        71928 => X"52",  -- 82
        71929 => X"5D",  -- 93
        71930 => X"76",  -- 118
        71931 => X"77",  -- 119
        71932 => X"64",  -- 100
        71933 => X"54",  -- 84
        71934 => X"79",  -- 121
        71935 => X"63",  -- 99
        71936 => X"74",  -- 116
        71937 => X"5B",  -- 91
        71938 => X"61",  -- 97
        71939 => X"6F",  -- 111
        71940 => X"6B",  -- 107
        71941 => X"74",  -- 116
        71942 => X"82",  -- 130
        71943 => X"7D",  -- 125
        71944 => X"59",  -- 89
        71945 => X"8C",  -- 140
        71946 => X"69",  -- 105
        71947 => X"52",  -- 82
        71948 => X"58",  -- 88
        71949 => X"8A",  -- 138
        71950 => X"7D",  -- 125
        71951 => X"86",  -- 134
        71952 => X"87",  -- 135
        71953 => X"8B",  -- 139
        71954 => X"8D",  -- 141
        71955 => X"89",  -- 137
        71956 => X"92",  -- 146
        71957 => X"90",  -- 144
        71958 => X"80",  -- 128
        71959 => X"8F",  -- 143
        71960 => X"98",  -- 152
        71961 => X"AA",  -- 170
        71962 => X"A4",  -- 164
        71963 => X"92",  -- 146
        71964 => X"8A",  -- 138
        71965 => X"7B",  -- 123
        71966 => X"6E",  -- 110
        71967 => X"69",  -- 105
        71968 => X"6A",  -- 106
        71969 => X"5C",  -- 92
        71970 => X"53",  -- 83
        71971 => X"57",  -- 87
        71972 => X"49",  -- 73
        71973 => X"4A",  -- 74
        71974 => X"3E",  -- 62
        71975 => X"4C",  -- 76
        71976 => X"7F",  -- 127
        71977 => X"8B",  -- 139
        71978 => X"7C",  -- 124
        71979 => X"7A",  -- 122
        71980 => X"8A",  -- 138
        71981 => X"7F",  -- 127
        71982 => X"56",  -- 86
        71983 => X"32",  -- 50
        71984 => X"3C",  -- 60
        71985 => X"4A",  -- 74
        71986 => X"67",  -- 103
        71987 => X"65",  -- 101
        71988 => X"7F",  -- 127
        71989 => X"75",  -- 117
        71990 => X"3B",  -- 59
        71991 => X"57",  -- 87
        71992 => X"5A",  -- 90
        71993 => X"54",  -- 84
        71994 => X"44",  -- 68
        71995 => X"38",  -- 56
        71996 => X"32",  -- 50
        71997 => X"2C",  -- 44
        71998 => X"3A",  -- 58
        71999 => X"56",  -- 86
        72000 => X"67",  -- 103
        72001 => X"66",  -- 102
        72002 => X"64",  -- 100
        72003 => X"61",  -- 97
        72004 => X"5E",  -- 94
        72005 => X"5F",  -- 95
        72006 => X"64",  -- 100
        72007 => X"69",  -- 105
        72008 => X"61",  -- 97
        72009 => X"59",  -- 89
        72010 => X"57",  -- 87
        72011 => X"5C",  -- 92
        72012 => X"5D",  -- 93
        72013 => X"58",  -- 88
        72014 => X"56",  -- 86
        72015 => X"59",  -- 89
        72016 => X"4E",  -- 78
        72017 => X"51",  -- 81
        72018 => X"57",  -- 87
        72019 => X"5F",  -- 95
        72020 => X"60",  -- 96
        72021 => X"5A",  -- 90
        72022 => X"53",  -- 83
        72023 => X"52",  -- 82
        72024 => X"54",  -- 84
        72025 => X"57",  -- 87
        72026 => X"4F",  -- 79
        72027 => X"3A",  -- 58
        72028 => X"4C",  -- 76
        72029 => X"69",  -- 105
        72030 => X"46",  -- 70
        72031 => X"47",  -- 71
        72032 => X"6B",  -- 107
        72033 => X"4F",  -- 79
        72034 => X"48",  -- 72
        72035 => X"45",  -- 69
        72036 => X"47",  -- 71
        72037 => X"49",  -- 73
        72038 => X"39",  -- 57
        72039 => X"33",  -- 51
        72040 => X"67",  -- 103
        72041 => X"45",  -- 69
        72042 => X"3A",  -- 58
        72043 => X"49",  -- 73
        72044 => X"49",  -- 73
        72045 => X"68",  -- 104
        72046 => X"52",  -- 82
        72047 => X"4C",  -- 76
        72048 => X"32",  -- 50
        72049 => X"2B",  -- 43
        72050 => X"24",  -- 36
        72051 => X"36",  -- 54
        72052 => X"32",  -- 50
        72053 => X"36",  -- 54
        72054 => X"26",  -- 38
        72055 => X"22",  -- 34
        72056 => X"21",  -- 33
        72057 => X"22",  -- 34
        72058 => X"24",  -- 36
        72059 => X"24",  -- 36
        72060 => X"1D",  -- 29
        72061 => X"17",  -- 23
        72062 => X"18",  -- 24
        72063 => X"1D",  -- 29
        72064 => X"2A",  -- 42
        72065 => X"22",  -- 34
        72066 => X"22",  -- 34
        72067 => X"2C",  -- 44
        72068 => X"2F",  -- 47
        72069 => X"27",  -- 39
        72070 => X"21",  -- 33
        72071 => X"21",  -- 33
        72072 => X"1E",  -- 30
        72073 => X"23",  -- 35
        72074 => X"28",  -- 40
        72075 => X"26",  -- 38
        72076 => X"20",  -- 32
        72077 => X"1C",  -- 28
        72078 => X"21",  -- 33
        72079 => X"26",  -- 38
        72080 => X"23",  -- 35
        72081 => X"18",  -- 24
        72082 => X"18",  -- 24
        72083 => X"1D",  -- 29
        72084 => X"1A",  -- 26
        72085 => X"1A",  -- 26
        72086 => X"1C",  -- 28
        72087 => X"19",  -- 25
        72088 => X"1A",  -- 26
        72089 => X"22",  -- 34
        72090 => X"28",  -- 40
        72091 => X"27",  -- 39
        72092 => X"23",  -- 35
        72093 => X"21",  -- 33
        72094 => X"1E",  -- 30
        72095 => X"1C",  -- 28
        72096 => X"1A",  -- 26
        72097 => X"1A",  -- 26
        72098 => X"1C",  -- 28
        72099 => X"1C",  -- 28
        72100 => X"17",  -- 23
        72101 => X"14",  -- 20
        72102 => X"18",  -- 24
        72103 => X"1E",  -- 30
        72104 => X"1C",  -- 28
        72105 => X"16",  -- 22
        72106 => X"17",  -- 23
        72107 => X"20",  -- 32
        72108 => X"24",  -- 36
        72109 => X"1E",  -- 30
        72110 => X"17",  -- 23
        72111 => X"17",  -- 23
        72112 => X"1C",  -- 28
        72113 => X"20",  -- 32
        72114 => X"2A",  -- 42
        72115 => X"2D",  -- 45
        72116 => X"25",  -- 37
        72117 => X"27",  -- 39
        72118 => X"30",  -- 48
        72119 => X"30",  -- 48
        72120 => X"34",  -- 52
        72121 => X"2F",  -- 47
        72122 => X"2D",  -- 45
        72123 => X"30",  -- 48
        72124 => X"30",  -- 48
        72125 => X"2C",  -- 44
        72126 => X"28",  -- 40
        72127 => X"28",  -- 40
        72128 => X"30",  -- 48
        72129 => X"29",  -- 41
        72130 => X"25",  -- 37
        72131 => X"29",  -- 41
        72132 => X"2E",  -- 46
        72133 => X"35",  -- 53
        72134 => X"3C",  -- 60
        72135 => X"44",  -- 68
        72136 => X"54",  -- 84
        72137 => X"4C",  -- 76
        72138 => X"3E",  -- 62
        72139 => X"34",  -- 52
        72140 => X"2F",  -- 47
        72141 => X"34",  -- 52
        72142 => X"3C",  -- 60
        72143 => X"41",  -- 65
        72144 => X"40",  -- 64
        72145 => X"59",  -- 89
        72146 => X"3E",  -- 62
        72147 => X"3C",  -- 60
        72148 => X"48",  -- 72
        72149 => X"3D",  -- 61
        72150 => X"43",  -- 67
        72151 => X"42",  -- 66
        72152 => X"49",  -- 73
        72153 => X"37",  -- 55
        72154 => X"3D",  -- 61
        72155 => X"47",  -- 71
        72156 => X"45",  -- 69
        72157 => X"4D",  -- 77
        72158 => X"4D",  -- 77
        72159 => X"36",  -- 54
        72160 => X"3C",  -- 60
        72161 => X"46",  -- 70
        72162 => X"49",  -- 73
        72163 => X"59",  -- 89
        72164 => X"61",  -- 97
        72165 => X"61",  -- 97
        72166 => X"6D",  -- 109
        72167 => X"6E",  -- 110
        72168 => X"66",  -- 102
        72169 => X"70",  -- 112
        72170 => X"78",  -- 120
        72171 => X"7B",  -- 123
        72172 => X"80",  -- 128
        72173 => X"87",  -- 135
        72174 => X"8B",  -- 139
        72175 => X"8D",  -- 141
        72176 => X"87",  -- 135
        72177 => X"82",  -- 130
        72178 => X"78",  -- 120
        72179 => X"70",  -- 112
        72180 => X"67",  -- 103
        72181 => X"5F",  -- 95
        72182 => X"57",  -- 87
        72183 => X"51",  -- 81
        72184 => X"64",  -- 100
        72185 => X"61",  -- 97
        72186 => X"5F",  -- 95
        72187 => X"60",  -- 96
        72188 => X"60",  -- 96
        72189 => X"61",  -- 97
        72190 => X"64",  -- 100
        72191 => X"67",  -- 103
        72192 => X"62",  -- 98
        72193 => X"64",  -- 100
        72194 => X"56",  -- 86
        72195 => X"50",  -- 80
        72196 => X"5D",  -- 93
        72197 => X"65",  -- 101
        72198 => X"62",  -- 98
        72199 => X"67",  -- 103
        72200 => X"61",  -- 97
        72201 => X"67",  -- 103
        72202 => X"66",  -- 102
        72203 => X"65",  -- 101
        72204 => X"66",  -- 102
        72205 => X"62",  -- 98
        72206 => X"5C",  -- 92
        72207 => X"5F",  -- 95
        72208 => X"5C",  -- 92
        72209 => X"5E",  -- 94
        72210 => X"5F",  -- 95
        72211 => X"5C",  -- 92
        72212 => X"56",  -- 86
        72213 => X"55",  -- 85
        72214 => X"5D",  -- 93
        72215 => X"67",  -- 103
        72216 => X"65",  -- 101
        72217 => X"6C",  -- 108
        72218 => X"55",  -- 85
        72219 => X"6C",  -- 108
        72220 => X"5E",  -- 94
        72221 => X"7B",  -- 123
        72222 => X"5A",  -- 90
        72223 => X"71",  -- 113
        72224 => X"6E",  -- 110
        72225 => X"58",  -- 88
        72226 => X"4E",  -- 78
        72227 => X"5C",  -- 92
        72228 => X"69",  -- 105
        72229 => X"64",  -- 100
        72230 => X"56",  -- 86
        72231 => X"50",  -- 80
        72232 => X"4C",  -- 76
        72233 => X"46",  -- 70
        72234 => X"4A",  -- 74
        72235 => X"5B",  -- 91
        72236 => X"64",  -- 100
        72237 => X"64",  -- 100
        72238 => X"66",  -- 102
        72239 => X"6C",  -- 108
        72240 => X"62",  -- 98
        72241 => X"5C",  -- 92
        72242 => X"66",  -- 102
        72243 => X"75",  -- 117
        72244 => X"75",  -- 117
        72245 => X"6D",  -- 109
        72246 => X"66",  -- 102
        72247 => X"62",  -- 98
        72248 => X"6E",  -- 110
        72249 => X"69",  -- 105
        72250 => X"64",  -- 100
        72251 => X"6A",  -- 106
        72252 => X"7D",  -- 125
        72253 => X"62",  -- 98
        72254 => X"66",  -- 102
        72255 => X"73",  -- 115
        72256 => X"77",  -- 119
        72257 => X"67",  -- 103
        72258 => X"77",  -- 119
        72259 => X"82",  -- 130
        72260 => X"6A",  -- 106
        72261 => X"59",  -- 89
        72262 => X"5E",  -- 94
        72263 => X"60",  -- 96
        72264 => X"61",  -- 97
        72265 => X"6B",  -- 107
        72266 => X"63",  -- 99
        72267 => X"80",  -- 128
        72268 => X"7B",  -- 123
        72269 => X"8B",  -- 139
        72270 => X"81",  -- 129
        72271 => X"96",  -- 150
        72272 => X"80",  -- 128
        72273 => X"80",  -- 128
        72274 => X"96",  -- 150
        72275 => X"81",  -- 129
        72276 => X"59",  -- 89
        72277 => X"6B",  -- 107
        72278 => X"8B",  -- 139
        72279 => X"96",  -- 150
        72280 => X"B4",  -- 180
        72281 => X"A3",  -- 163
        72282 => X"9C",  -- 156
        72283 => X"87",  -- 135
        72284 => X"59",  -- 89
        72285 => X"61",  -- 97
        72286 => X"51",  -- 81
        72287 => X"5D",  -- 93
        72288 => X"60",  -- 96
        72289 => X"64",  -- 100
        72290 => X"5B",  -- 91
        72291 => X"4C",  -- 76
        72292 => X"3E",  -- 62
        72293 => X"5F",  -- 95
        72294 => X"59",  -- 89
        72295 => X"45",  -- 69
        72296 => X"69",  -- 105
        72297 => X"80",  -- 128
        72298 => X"75",  -- 117
        72299 => X"65",  -- 101
        72300 => X"75",  -- 117
        72301 => X"7A",  -- 122
        72302 => X"54",  -- 84
        72303 => X"23",  -- 35
        72304 => X"30",  -- 48
        72305 => X"37",  -- 55
        72306 => X"57",  -- 87
        72307 => X"61",  -- 97
        72308 => X"56",  -- 86
        72309 => X"4E",  -- 78
        72310 => X"4A",  -- 74
        72311 => X"52",  -- 82
        72312 => X"52",  -- 82
        72313 => X"52",  -- 82
        72314 => X"4C",  -- 76
        72315 => X"47",  -- 71
        72316 => X"42",  -- 66
        72317 => X"37",  -- 55
        72318 => X"3A",  -- 58
        72319 => X"4C",  -- 76
        72320 => X"6C",  -- 108
        72321 => X"6F",  -- 111
        72322 => X"68",  -- 104
        72323 => X"5B",  -- 91
        72324 => X"5B",  -- 91
        72325 => X"66",  -- 102
        72326 => X"68",  -- 104
        72327 => X"60",  -- 96
        72328 => X"5B",  -- 91
        72329 => X"5B",  -- 91
        72330 => X"58",  -- 88
        72331 => X"54",  -- 84
        72332 => X"50",  -- 80
        72333 => X"53",  -- 83
        72334 => X"5A",  -- 90
        72335 => X"60",  -- 96
        72336 => X"5B",  -- 91
        72337 => X"56",  -- 86
        72338 => X"59",  -- 89
        72339 => X"60",  -- 96
        72340 => X"5B",  -- 91
        72341 => X"4E",  -- 78
        72342 => X"49",  -- 73
        72343 => X"4B",  -- 75
        72344 => X"46",  -- 70
        72345 => X"4F",  -- 79
        72346 => X"56",  -- 86
        72347 => X"3F",  -- 63
        72348 => X"65",  -- 101
        72349 => X"52",  -- 82
        72350 => X"47",  -- 71
        72351 => X"3E",  -- 62
        72352 => X"63",  -- 99
        72353 => X"53",  -- 83
        72354 => X"52",  -- 82
        72355 => X"4C",  -- 76
        72356 => X"4C",  -- 76
        72357 => X"4A",  -- 74
        72358 => X"38",  -- 56
        72359 => X"34",  -- 52
        72360 => X"6E",  -- 110
        72361 => X"37",  -- 55
        72362 => X"3C",  -- 60
        72363 => X"4A",  -- 74
        72364 => X"4B",  -- 75
        72365 => X"7A",  -- 122
        72366 => X"4D",  -- 77
        72367 => X"65",  -- 101
        72368 => X"31",  -- 49
        72369 => X"28",  -- 40
        72370 => X"24",  -- 36
        72371 => X"35",  -- 53
        72372 => X"37",  -- 55
        72373 => X"40",  -- 64
        72374 => X"35",  -- 53
        72375 => X"29",  -- 41
        72376 => X"23",  -- 35
        72377 => X"23",  -- 35
        72378 => X"25",  -- 37
        72379 => X"24",  -- 36
        72380 => X"1F",  -- 31
        72381 => X"1A",  -- 26
        72382 => X"1C",  -- 28
        72383 => X"21",  -- 33
        72384 => X"2B",  -- 43
        72385 => X"22",  -- 34
        72386 => X"1E",  -- 30
        72387 => X"25",  -- 37
        72388 => X"2E",  -- 46
        72389 => X"2E",  -- 46
        72390 => X"27",  -- 39
        72391 => X"22",  -- 34
        72392 => X"23",  -- 35
        72393 => X"28",  -- 40
        72394 => X"2A",  -- 42
        72395 => X"25",  -- 37
        72396 => X"1D",  -- 29
        72397 => X"18",  -- 24
        72398 => X"1B",  -- 27
        72399 => X"1F",  -- 31
        72400 => X"25",  -- 37
        72401 => X"20",  -- 32
        72402 => X"24",  -- 36
        72403 => X"24",  -- 36
        72404 => X"1B",  -- 27
        72405 => X"19",  -- 25
        72406 => X"1F",  -- 31
        72407 => X"1F",  -- 31
        72408 => X"1D",  -- 29
        72409 => X"25",  -- 37
        72410 => X"2B",  -- 43
        72411 => X"27",  -- 39
        72412 => X"21",  -- 33
        72413 => X"1D",  -- 29
        72414 => X"1C",  -- 28
        72415 => X"19",  -- 25
        72416 => X"19",  -- 25
        72417 => X"19",  -- 25
        72418 => X"1B",  -- 27
        72419 => X"1C",  -- 28
        72420 => X"18",  -- 24
        72421 => X"16",  -- 22
        72422 => X"1B",  -- 27
        72423 => X"22",  -- 34
        72424 => X"19",  -- 25
        72425 => X"15",  -- 21
        72426 => X"17",  -- 23
        72427 => X"20",  -- 32
        72428 => X"23",  -- 35
        72429 => X"1C",  -- 28
        72430 => X"15",  -- 21
        72431 => X"15",  -- 21
        72432 => X"14",  -- 20
        72433 => X"1C",  -- 28
        72434 => X"29",  -- 41
        72435 => X"2B",  -- 43
        72436 => X"25",  -- 37
        72437 => X"29",  -- 41
        72438 => X"2E",  -- 46
        72439 => X"28",  -- 40
        72440 => X"25",  -- 37
        72441 => X"25",  -- 37
        72442 => X"29",  -- 41
        72443 => X"31",  -- 49
        72444 => X"36",  -- 54
        72445 => X"34",  -- 52
        72446 => X"30",  -- 48
        72447 => X"2D",  -- 45
        72448 => X"28",  -- 40
        72449 => X"24",  -- 36
        72450 => X"22",  -- 34
        72451 => X"23",  -- 35
        72452 => X"23",  -- 35
        72453 => X"25",  -- 37
        72454 => X"2D",  -- 45
        72455 => X"34",  -- 52
        72456 => X"3F",  -- 63
        72457 => X"40",  -- 64
        72458 => X"40",  -- 64
        72459 => X"3F",  -- 63
        72460 => X"3D",  -- 61
        72461 => X"3C",  -- 60
        72462 => X"3F",  -- 63
        72463 => X"42",  -- 66
        72464 => X"38",  -- 56
        72465 => X"4E",  -- 78
        72466 => X"4C",  -- 76
        72467 => X"42",  -- 66
        72468 => X"44",  -- 68
        72469 => X"41",  -- 65
        72470 => X"3C",  -- 60
        72471 => X"45",  -- 69
        72472 => X"41",  -- 65
        72473 => X"39",  -- 57
        72474 => X"45",  -- 69
        72475 => X"52",  -- 82
        72476 => X"49",  -- 73
        72477 => X"47",  -- 71
        72478 => X"4D",  -- 77
        72479 => X"46",  -- 70
        72480 => X"3F",  -- 63
        72481 => X"52",  -- 82
        72482 => X"5B",  -- 91
        72483 => X"69",  -- 105
        72484 => X"6D",  -- 109
        72485 => X"6E",  -- 110
        72486 => X"7A",  -- 122
        72487 => X"7A",  -- 122
        72488 => X"7B",  -- 123
        72489 => X"7D",  -- 125
        72490 => X"80",  -- 128
        72491 => X"85",  -- 133
        72492 => X"8D",  -- 141
        72493 => X"96",  -- 150
        72494 => X"9C",  -- 156
        72495 => X"9D",  -- 157
        72496 => X"9C",  -- 156
        72497 => X"9D",  -- 157
        72498 => X"93",  -- 147
        72499 => X"7F",  -- 127
        72500 => X"6F",  -- 111
        72501 => X"66",  -- 102
        72502 => X"5D",  -- 93
        72503 => X"53",  -- 83
        72504 => X"64",  -- 100
        72505 => X"60",  -- 96
        72506 => X"61",  -- 97
        72507 => X"5D",  -- 93
        72508 => X"55",  -- 85
        72509 => X"61",  -- 97
        72510 => X"6B",  -- 107
        72511 => X"61",  -- 97
        72512 => X"5F",  -- 95
        72513 => X"60",  -- 96
        72514 => X"55",  -- 85
        72515 => X"50",  -- 80
        72516 => X"5C",  -- 92
        72517 => X"61",  -- 97
        72518 => X"5D",  -- 93
        72519 => X"5F",  -- 95
        72520 => X"5D",  -- 93
        72521 => X"60",  -- 96
        72522 => X"62",  -- 98
        72523 => X"66",  -- 102
        72524 => X"6A",  -- 106
        72525 => X"60",  -- 96
        72526 => X"5B",  -- 91
        72527 => X"61",  -- 97
        72528 => X"6F",  -- 111
        72529 => X"6F",  -- 111
        72530 => X"72",  -- 114
        72531 => X"71",  -- 113
        72532 => X"6C",  -- 108
        72533 => X"66",  -- 102
        72534 => X"6D",  -- 109
        72535 => X"76",  -- 118
        72536 => X"63",  -- 99
        72537 => X"69",  -- 105
        72538 => X"59",  -- 89
        72539 => X"6D",  -- 109
        72540 => X"5C",  -- 92
        72541 => X"74",  -- 116
        72542 => X"58",  -- 88
        72543 => X"6D",  -- 109
        72544 => X"4D",  -- 77
        72545 => X"3B",  -- 59
        72546 => X"36",  -- 54
        72547 => X"48",  -- 72
        72548 => X"5A",  -- 90
        72549 => X"59",  -- 89
        72550 => X"4E",  -- 78
        72551 => X"46",  -- 70
        72552 => X"48",  -- 72
        72553 => X"42",  -- 66
        72554 => X"4C",  -- 76
        72555 => X"5E",  -- 94
        72556 => X"64",  -- 100
        72557 => X"5B",  -- 91
        72558 => X"5B",  -- 91
        72559 => X"68",  -- 104
        72560 => X"57",  -- 87
        72561 => X"5A",  -- 90
        72562 => X"65",  -- 101
        72563 => X"77",  -- 119
        72564 => X"84",  -- 132
        72565 => X"83",  -- 131
        72566 => X"86",  -- 134
        72567 => X"94",  -- 148
        72568 => X"74",  -- 116
        72569 => X"76",  -- 118
        72570 => X"73",  -- 115
        72571 => X"5E",  -- 94
        72572 => X"69",  -- 105
        72573 => X"6B",  -- 107
        72574 => X"6B",  -- 107
        72575 => X"77",  -- 119
        72576 => X"53",  -- 83
        72577 => X"59",  -- 89
        72578 => X"70",  -- 112
        72579 => X"75",  -- 117
        72580 => X"5F",  -- 95
        72581 => X"5B",  -- 91
        72582 => X"6D",  -- 109
        72583 => X"78",  -- 120
        72584 => X"59",  -- 89
        72585 => X"4E",  -- 78
        72586 => X"51",  -- 81
        72587 => X"74",  -- 116
        72588 => X"66",  -- 102
        72589 => X"74",  -- 116
        72590 => X"74",  -- 116
        72591 => X"79",  -- 121
        72592 => X"77",  -- 119
        72593 => X"7A",  -- 122
        72594 => X"74",  -- 116
        72595 => X"5A",  -- 90
        72596 => X"53",  -- 83
        72597 => X"69",  -- 105
        72598 => X"84",  -- 132
        72599 => X"A8",  -- 168
        72600 => X"98",  -- 152
        72601 => X"7B",  -- 123
        72602 => X"8E",  -- 142
        72603 => X"8F",  -- 143
        72604 => X"4E",  -- 78
        72605 => X"52",  -- 82
        72606 => X"36",  -- 54
        72607 => X"43",  -- 67
        72608 => X"56",  -- 86
        72609 => X"51",  -- 81
        72610 => X"49",  -- 73
        72611 => X"48",  -- 72
        72612 => X"3A",  -- 58
        72613 => X"5F",  -- 95
        72614 => X"65",  -- 101
        72615 => X"4F",  -- 79
        72616 => X"4D",  -- 77
        72617 => X"63",  -- 99
        72618 => X"62",  -- 98
        72619 => X"58",  -- 88
        72620 => X"68",  -- 104
        72621 => X"78",  -- 120
        72622 => X"67",  -- 103
        72623 => X"4D",  -- 77
        72624 => X"54",  -- 84
        72625 => X"4B",  -- 75
        72626 => X"48",  -- 72
        72627 => X"5F",  -- 95
        72628 => X"64",  -- 100
        72629 => X"61",  -- 97
        72630 => X"68",  -- 104
        72631 => X"58",  -- 88
        72632 => X"46",  -- 70
        72633 => X"4D",  -- 77
        72634 => X"4F",  -- 79
        72635 => X"50",  -- 80
        72636 => X"50",  -- 80
        72637 => X"46",  -- 70
        72638 => X"42",  -- 66
        72639 => X"4D",  -- 77
        72640 => X"66",  -- 102
        72641 => X"6C",  -- 108
        72642 => X"6A",  -- 106
        72643 => X"61",  -- 97
        72644 => X"60",  -- 96
        72645 => X"65",  -- 101
        72646 => X"63",  -- 99
        72647 => X"58",  -- 88
        72648 => X"5A",  -- 90
        72649 => X"5D",  -- 93
        72650 => X"5A",  -- 90
        72651 => X"4F",  -- 79
        72652 => X"49",  -- 73
        72653 => X"50",  -- 80
        72654 => X"58",  -- 88
        72655 => X"5B",  -- 91
        72656 => X"5C",  -- 92
        72657 => X"56",  -- 86
        72658 => X"57",  -- 87
        72659 => X"5C",  -- 92
        72660 => X"55",  -- 85
        72661 => X"45",  -- 69
        72662 => X"42",  -- 66
        72663 => X"4A",  -- 74
        72664 => X"49",  -- 73
        72665 => X"4B",  -- 75
        72666 => X"53",  -- 83
        72667 => X"5B",  -- 91
        72668 => X"7D",  -- 125
        72669 => X"42",  -- 66
        72670 => X"3D",  -- 61
        72671 => X"39",  -- 57
        72672 => X"4C",  -- 76
        72673 => X"4F",  -- 79
        72674 => X"5B",  -- 91
        72675 => X"52",  -- 82
        72676 => X"4A",  -- 74
        72677 => X"44",  -- 68
        72678 => X"39",  -- 57
        72679 => X"45",  -- 69
        72680 => X"65",  -- 101
        72681 => X"34",  -- 52
        72682 => X"40",  -- 64
        72683 => X"58",  -- 88
        72684 => X"5A",  -- 90
        72685 => X"80",  -- 128
        72686 => X"4D",  -- 77
        72687 => X"71",  -- 113
        72688 => X"42",  -- 66
        72689 => X"31",  -- 49
        72690 => X"2B",  -- 43
        72691 => X"31",  -- 49
        72692 => X"32",  -- 50
        72693 => X"3F",  -- 63
        72694 => X"42",  -- 66
        72695 => X"36",  -- 54
        72696 => X"21",  -- 33
        72697 => X"22",  -- 34
        72698 => X"25",  -- 37
        72699 => X"28",  -- 40
        72700 => X"25",  -- 37
        72701 => X"21",  -- 33
        72702 => X"22",  -- 34
        72703 => X"27",  -- 39
        72704 => X"24",  -- 36
        72705 => X"2D",  -- 45
        72706 => X"2B",  -- 43
        72707 => X"24",  -- 36
        72708 => X"2C",  -- 44
        72709 => X"39",  -- 57
        72710 => X"30",  -- 48
        72711 => X"1A",  -- 26
        72712 => X"21",  -- 33
        72713 => X"2C",  -- 44
        72714 => X"31",  -- 49
        72715 => X"2A",  -- 42
        72716 => X"1D",  -- 29
        72717 => X"16",  -- 22
        72718 => X"18",  -- 24
        72719 => X"1C",  -- 28
        72720 => X"21",  -- 33
        72721 => X"25",  -- 37
        72722 => X"31",  -- 49
        72723 => X"35",  -- 53
        72724 => X"2A",  -- 42
        72725 => X"22",  -- 34
        72726 => X"20",  -- 32
        72727 => X"1A",  -- 26
        72728 => X"19",  -- 25
        72729 => X"21",  -- 33
        72730 => X"27",  -- 39
        72731 => X"24",  -- 36
        72732 => X"1D",  -- 29
        72733 => X"1B",  -- 27
        72734 => X"1C",  -- 28
        72735 => X"1C",  -- 28
        72736 => X"19",  -- 25
        72737 => X"18",  -- 24
        72738 => X"1A",  -- 26
        72739 => X"19",  -- 25
        72740 => X"15",  -- 21
        72741 => X"12",  -- 18
        72742 => X"16",  -- 22
        72743 => X"1D",  -- 29
        72744 => X"1A",  -- 26
        72745 => X"16",  -- 22
        72746 => X"17",  -- 23
        72747 => X"1D",  -- 29
        72748 => X"1E",  -- 30
        72749 => X"17",  -- 23
        72750 => X"12",  -- 18
        72751 => X"14",  -- 20
        72752 => X"12",  -- 18
        72753 => X"1D",  -- 29
        72754 => X"2B",  -- 43
        72755 => X"2C",  -- 44
        72756 => X"27",  -- 39
        72757 => X"2C",  -- 44
        72758 => X"30",  -- 48
        72759 => X"27",  -- 39
        72760 => X"1D",  -- 29
        72761 => X"1F",  -- 31
        72762 => X"25",  -- 37
        72763 => X"2E",  -- 46
        72764 => X"35",  -- 53
        72765 => X"37",  -- 55
        72766 => X"34",  -- 52
        72767 => X"30",  -- 48
        72768 => X"29",  -- 41
        72769 => X"28",  -- 40
        72770 => X"25",  -- 37
        72771 => X"21",  -- 33
        72772 => X"1D",  -- 29
        72773 => X"1E",  -- 30
        72774 => X"26",  -- 38
        72775 => X"2D",  -- 45
        72776 => X"2D",  -- 45
        72777 => X"35",  -- 53
        72778 => X"3E",  -- 62
        72779 => X"40",  -- 64
        72780 => X"3F",  -- 63
        72781 => X"3C",  -- 60
        72782 => X"3B",  -- 59
        72783 => X"3D",  -- 61
        72784 => X"2F",  -- 47
        72785 => X"41",  -- 65
        72786 => X"55",  -- 85
        72787 => X"49",  -- 73
        72788 => X"47",  -- 71
        72789 => X"44",  -- 68
        72790 => X"30",  -- 48
        72791 => X"37",  -- 55
        72792 => X"32",  -- 50
        72793 => X"36",  -- 54
        72794 => X"48",  -- 72
        72795 => X"52",  -- 82
        72796 => X"49",  -- 73
        72797 => X"4C",  -- 76
        72798 => X"58",  -- 88
        72799 => X"5A",  -- 90
        72800 => X"53",  -- 83
        72801 => X"66",  -- 102
        72802 => X"6C",  -- 108
        72803 => X"75",  -- 117
        72804 => X"75",  -- 117
        72805 => X"74",  -- 116
        72806 => X"7E",  -- 126
        72807 => X"7B",  -- 123
        72808 => X"7D",  -- 125
        72809 => X"7E",  -- 126
        72810 => X"7F",  -- 127
        72811 => X"82",  -- 130
        72812 => X"86",  -- 134
        72813 => X"8E",  -- 142
        72814 => X"94",  -- 148
        72815 => X"97",  -- 151
        72816 => X"99",  -- 153
        72817 => X"A2",  -- 162
        72818 => X"9D",  -- 157
        72819 => X"8C",  -- 140
        72820 => X"7B",  -- 123
        72821 => X"6F",  -- 111
        72822 => X"5D",  -- 93
        72823 => X"4D",  -- 77
        72824 => X"53",  -- 83
        72825 => X"55",  -- 85
        72826 => X"61",  -- 97
        72827 => X"58",  -- 88
        72828 => X"45",  -- 69
        72829 => X"51",  -- 81
        72830 => X"61",  -- 97
        72831 => X"52",  -- 82
        72832 => X"59",  -- 89
        72833 => X"5A",  -- 90
        72834 => X"58",  -- 88
        72835 => X"56",  -- 86
        72836 => X"5A",  -- 90
        72837 => X"5B",  -- 91
        72838 => X"59",  -- 89
        72839 => X"5A",  -- 90
        72840 => X"5B",  -- 91
        72841 => X"5B",  -- 91
        72842 => X"5D",  -- 93
        72843 => X"65",  -- 101
        72844 => X"6C",  -- 108
        72845 => X"61",  -- 97
        72846 => X"5D",  -- 93
        72847 => X"69",  -- 105
        72848 => X"73",  -- 115
        72849 => X"6E",  -- 110
        72850 => X"70",  -- 112
        72851 => X"76",  -- 118
        72852 => X"75",  -- 117
        72853 => X"6B",  -- 107
        72854 => X"66",  -- 102
        72855 => X"68",  -- 104
        72856 => X"4C",  -- 76
        72857 => X"45",  -- 69
        72858 => X"4A",  -- 74
        72859 => X"49",  -- 73
        72860 => X"4E",  -- 78
        72861 => X"4F",  -- 79
        72862 => X"43",  -- 67
        72863 => X"46",  -- 70
        72864 => X"30",  -- 48
        72865 => X"31",  -- 49
        72866 => X"3B",  -- 59
        72867 => X"49",  -- 73
        72868 => X"52",  -- 82
        72869 => X"4D",  -- 77
        72870 => X"47",  -- 71
        72871 => X"45",  -- 69
        72872 => X"47",  -- 71
        72873 => X"44",  -- 68
        72874 => X"4A",  -- 74
        72875 => X"57",  -- 87
        72876 => X"5C",  -- 92
        72877 => X"56",  -- 86
        72878 => X"57",  -- 87
        72879 => X"5F",  -- 95
        72880 => X"65",  -- 101
        72881 => X"69",  -- 105
        72882 => X"64",  -- 100
        72883 => X"66",  -- 102
        72884 => X"78",  -- 120
        72885 => X"7C",  -- 124
        72886 => X"79",  -- 121
        72887 => X"83",  -- 131
        72888 => X"78",  -- 120
        72889 => X"6A",  -- 106
        72890 => X"7B",  -- 123
        72891 => X"5E",  -- 94
        72892 => X"48",  -- 72
        72893 => X"66",  -- 102
        72894 => X"76",  -- 118
        72895 => X"6C",  -- 108
        72896 => X"64",  -- 100
        72897 => X"72",  -- 114
        72898 => X"7B",  -- 123
        72899 => X"6B",  -- 107
        72900 => X"54",  -- 84
        72901 => X"5A",  -- 90
        72902 => X"68",  -- 104
        72903 => X"64",  -- 100
        72904 => X"6A",  -- 106
        72905 => X"5A",  -- 90
        72906 => X"49",  -- 73
        72907 => X"54",  -- 84
        72908 => X"51",  -- 81
        72909 => X"6D",  -- 109
        72910 => X"74",  -- 116
        72911 => X"76",  -- 118
        72912 => X"8B",  -- 139
        72913 => X"79",  -- 121
        72914 => X"5E",  -- 94
        72915 => X"4D",  -- 77
        72916 => X"60",  -- 96
        72917 => X"6A",  -- 106
        72918 => X"6D",  -- 109
        72919 => X"92",  -- 146
        72920 => X"94",  -- 148
        72921 => X"7A",  -- 122
        72922 => X"88",  -- 136
        72923 => X"91",  -- 145
        72924 => X"62",  -- 98
        72925 => X"4D",  -- 77
        72926 => X"39",  -- 57
        72927 => X"47",  -- 71
        72928 => X"4D",  -- 77
        72929 => X"3F",  -- 63
        72930 => X"3B",  -- 59
        72931 => X"4A",  -- 74
        72932 => X"3B",  -- 59
        72933 => X"59",  -- 89
        72934 => X"6E",  -- 110
        72935 => X"5F",  -- 95
        72936 => X"36",  -- 54
        72937 => X"3B",  -- 59
        72938 => X"50",  -- 80
        72939 => X"66",  -- 102
        72940 => X"76",  -- 118
        72941 => X"76",  -- 118
        72942 => X"70",  -- 112
        72943 => X"79",  -- 121
        72944 => X"54",  -- 84
        72945 => X"67",  -- 103
        72946 => X"5B",  -- 91
        72947 => X"60",  -- 96
        72948 => X"6E",  -- 110
        72949 => X"5E",  -- 94
        72950 => X"5A",  -- 90
        72951 => X"6B",  -- 107
        72952 => X"4F",  -- 79
        72953 => X"56",  -- 86
        72954 => X"54",  -- 84
        72955 => X"51",  -- 81
        72956 => X"52",  -- 82
        72957 => X"4C",  -- 76
        72958 => X"48",  -- 72
        72959 => X"4F",  -- 79
        72960 => X"5F",  -- 95
        72961 => X"61",  -- 97
        72962 => X"66",  -- 102
        72963 => X"68",  -- 104
        72964 => X"63",  -- 99
        72965 => X"5C",  -- 92
        72966 => X"59",  -- 89
        72967 => X"5B",  -- 91
        72968 => X"5E",  -- 94
        72969 => X"62",  -- 98
        72970 => X"5E",  -- 94
        72971 => X"54",  -- 84
        72972 => X"51",  -- 81
        72973 => X"58",  -- 88
        72974 => X"5B",  -- 91
        72975 => X"58",  -- 88
        72976 => X"54",  -- 84
        72977 => X"51",  -- 81
        72978 => X"54",  -- 84
        72979 => X"58",  -- 88
        72980 => X"51",  -- 81
        72981 => X"46",  -- 70
        72982 => X"46",  -- 70
        72983 => X"4F",  -- 79
        72984 => X"59",  -- 89
        72985 => X"5A",  -- 90
        72986 => X"53",  -- 83
        72987 => X"72",  -- 114
        72988 => X"76",  -- 118
        72989 => X"44",  -- 68
        72990 => X"3A",  -- 58
        72991 => X"36",  -- 54
        72992 => X"4A",  -- 74
        72993 => X"51",  -- 81
        72994 => X"5D",  -- 93
        72995 => X"54",  -- 84
        72996 => X"4D",  -- 77
        72997 => X"44",  -- 68
        72998 => X"3D",  -- 61
        72999 => X"54",  -- 84
        73000 => X"57",  -- 87
        73001 => X"3F",  -- 63
        73002 => X"48",  -- 72
        73003 => X"6A",  -- 106
        73004 => X"68",  -- 104
        73005 => X"71",  -- 113
        73006 => X"47",  -- 71
        73007 => X"5F",  -- 95
        73008 => X"4E",  -- 78
        73009 => X"37",  -- 55
        73010 => X"33",  -- 51
        73011 => X"30",  -- 48
        73012 => X"2B",  -- 43
        73013 => X"34",  -- 52
        73014 => X"41",  -- 65
        73015 => X"37",  -- 55
        73016 => X"20",  -- 32
        73017 => X"21",  -- 33
        73018 => X"25",  -- 37
        73019 => X"29",  -- 41
        73020 => X"28",  -- 40
        73021 => X"24",  -- 36
        73022 => X"24",  -- 36
        73023 => X"27",  -- 39
        73024 => X"26",  -- 38
        73025 => X"34",  -- 52
        73026 => X"39",  -- 57
        73027 => X"33",  -- 51
        73028 => X"34",  -- 52
        73029 => X"39",  -- 57
        73030 => X"2E",  -- 46
        73031 => X"1A",  -- 26
        73032 => X"21",  -- 33
        73033 => X"34",  -- 52
        73034 => X"41",  -- 65
        73035 => X"39",  -- 57
        73036 => X"26",  -- 38
        73037 => X"1C",  -- 28
        73038 => X"1C",  -- 28
        73039 => X"20",  -- 32
        73040 => X"1C",  -- 28
        73041 => X"23",  -- 35
        73042 => X"33",  -- 51
        73043 => X"3C",  -- 60
        73044 => X"36",  -- 54
        73045 => X"2F",  -- 47
        73046 => X"27",  -- 39
        73047 => X"1B",  -- 27
        73048 => X"1B",  -- 27
        73049 => X"23",  -- 35
        73050 => X"28",  -- 40
        73051 => X"25",  -- 37
        73052 => X"20",  -- 32
        73053 => X"1F",  -- 31
        73054 => X"21",  -- 33
        73055 => X"21",  -- 33
        73056 => X"1B",  -- 27
        73057 => X"1A",  -- 26
        73058 => X"1A",  -- 26
        73059 => X"19",  -- 25
        73060 => X"14",  -- 20
        73061 => X"12",  -- 18
        73062 => X"16",  -- 22
        73063 => X"1E",  -- 30
        73064 => X"22",  -- 34
        73065 => X"1D",  -- 29
        73066 => X"1B",  -- 27
        73067 => X"1E",  -- 30
        73068 => X"1B",  -- 27
        73069 => X"14",  -- 20
        73070 => X"13",  -- 19
        73071 => X"18",  -- 24
        73072 => X"17",  -- 23
        73073 => X"1F",  -- 31
        73074 => X"2C",  -- 44
        73075 => X"30",  -- 48
        73076 => X"2D",  -- 45
        73077 => X"32",  -- 50
        73078 => X"35",  -- 53
        73079 => X"2D",  -- 45
        73080 => X"29",  -- 41
        73081 => X"29",  -- 41
        73082 => X"2A",  -- 42
        73083 => X"2C",  -- 44
        73084 => X"2F",  -- 47
        73085 => X"30",  -- 48
        73086 => X"2C",  -- 44
        73087 => X"28",  -- 40
        73088 => X"2A",  -- 42
        73089 => X"2B",  -- 43
        73090 => X"2B",  -- 43
        73091 => X"27",  -- 39
        73092 => X"24",  -- 36
        73093 => X"28",  -- 40
        73094 => X"31",  -- 49
        73095 => X"38",  -- 56
        73096 => X"30",  -- 48
        73097 => X"33",  -- 51
        73098 => X"36",  -- 54
        73099 => X"34",  -- 52
        73100 => X"31",  -- 49
        73101 => X"2F",  -- 47
        73102 => X"32",  -- 50
        73103 => X"36",  -- 54
        73104 => X"30",  -- 48
        73105 => X"36",  -- 54
        73106 => X"4C",  -- 76
        73107 => X"3C",  -- 60
        73108 => X"37",  -- 55
        73109 => X"3C",  -- 60
        73110 => X"27",  -- 39
        73111 => X"2C",  -- 44
        73112 => X"35",  -- 53
        73113 => X"3A",  -- 58
        73114 => X"44",  -- 68
        73115 => X"4B",  -- 75
        73116 => X"55",  -- 85
        73117 => X"66",  -- 102
        73118 => X"6C",  -- 108
        73119 => X"63",  -- 99
        73120 => X"6A",  -- 106
        73121 => X"74",  -- 116
        73122 => X"72",  -- 114
        73123 => X"78",  -- 120
        73124 => X"78",  -- 120
        73125 => X"75",  -- 117
        73126 => X"7D",  -- 125
        73127 => X"76",  -- 118
        73128 => X"75",  -- 117
        73129 => X"75",  -- 117
        73130 => X"76",  -- 118
        73131 => X"75",  -- 117
        73132 => X"73",  -- 115
        73133 => X"74",  -- 116
        73134 => X"7A",  -- 122
        73135 => X"81",  -- 129
        73136 => X"85",  -- 133
        73137 => X"90",  -- 144
        73138 => X"95",  -- 149
        73139 => X"90",  -- 144
        73140 => X"89",  -- 137
        73141 => X"7D",  -- 125
        73142 => X"63",  -- 99
        73143 => X"4B",  -- 75
        73144 => X"3A",  -- 58
        73145 => X"43",  -- 67
        73146 => X"5B",  -- 91
        73147 => X"5A",  -- 90
        73148 => X"40",  -- 64
        73149 => X"46",  -- 70
        73150 => X"56",  -- 86
        73151 => X"4E",  -- 78
        73152 => X"4D",  -- 77
        73153 => X"51",  -- 81
        73154 => X"59",  -- 89
        73155 => X"5B",  -- 91
        73156 => X"57",  -- 87
        73157 => X"53",  -- 83
        73158 => X"55",  -- 85
        73159 => X"56",  -- 86
        73160 => X"5D",  -- 93
        73161 => X"5C",  -- 92
        73162 => X"5C",  -- 92
        73163 => X"64",  -- 100
        73164 => X"68",  -- 104
        73165 => X"60",  -- 96
        73166 => X"5E",  -- 94
        73167 => X"6B",  -- 107
        73168 => X"6F",  -- 111
        73169 => X"6C",  -- 108
        73170 => X"6E",  -- 110
        73171 => X"70",  -- 112
        73172 => X"68",  -- 104
        73173 => X"5B",  -- 91
        73174 => X"55",  -- 85
        73175 => X"58",  -- 88
        73176 => X"48",  -- 72
        73177 => X"3B",  -- 59
        73178 => X"45",  -- 69
        73179 => X"46",  -- 70
        73180 => X"50",  -- 80
        73181 => X"4F",  -- 79
        73182 => X"44",  -- 68
        73183 => X"3F",  -- 63
        73184 => X"37",  -- 55
        73185 => X"40",  -- 64
        73186 => X"4B",  -- 75
        73187 => X"52",  -- 82
        73188 => X"4F",  -- 79
        73189 => X"49",  -- 73
        73190 => X"45",  -- 69
        73191 => X"45",  -- 69
        73192 => X"44",  -- 68
        73193 => X"48",  -- 72
        73194 => X"4B",  -- 75
        73195 => X"4F",  -- 79
        73196 => X"56",  -- 86
        73197 => X"57",  -- 87
        73198 => X"54",  -- 84
        73199 => X"4F",  -- 79
        73200 => X"55",  -- 85
        73201 => X"5F",  -- 95
        73202 => X"54",  -- 84
        73203 => X"49",  -- 73
        73204 => X"55",  -- 85
        73205 => X"62",  -- 98
        73206 => X"65",  -- 101
        73207 => X"6C",  -- 108
        73208 => X"7E",  -- 126
        73209 => X"59",  -- 89
        73210 => X"63",  -- 99
        73211 => X"5F",  -- 95
        73212 => X"4D",  -- 77
        73213 => X"62",  -- 98
        73214 => X"67",  -- 103
        73215 => X"67",  -- 103
        73216 => X"56",  -- 86
        73217 => X"5E",  -- 94
        73218 => X"68",  -- 104
        73219 => X"6D",  -- 109
        73220 => X"6F",  -- 111
        73221 => X"79",  -- 121
        73222 => X"7E",  -- 126
        73223 => X"78",  -- 120
        73224 => X"77",  -- 119
        73225 => X"63",  -- 99
        73226 => X"42",  -- 66
        73227 => X"49",  -- 73
        73228 => X"5C",  -- 92
        73229 => X"72",  -- 114
        73230 => X"76",  -- 118
        73231 => X"84",  -- 132
        73232 => X"66",  -- 102
        73233 => X"4A",  -- 74
        73234 => X"53",  -- 83
        73235 => X"57",  -- 87
        73236 => X"5A",  -- 90
        73237 => X"7C",  -- 124
        73238 => X"9B",  -- 155
        73239 => X"A5",  -- 165
        73240 => X"A5",  -- 165
        73241 => X"A1",  -- 161
        73242 => X"9C",  -- 156
        73243 => X"A2",  -- 162
        73244 => X"95",  -- 149
        73245 => X"53",  -- 83
        73246 => X"48",  -- 72
        73247 => X"45",  -- 69
        73248 => X"49",  -- 73
        73249 => X"4E",  -- 78
        73250 => X"4A",  -- 74
        73251 => X"52",  -- 82
        73252 => X"3B",  -- 59
        73253 => X"5A",  -- 90
        73254 => X"78",  -- 120
        73255 => X"64",  -- 100
        73256 => X"32",  -- 50
        73257 => X"23",  -- 35
        73258 => X"43",  -- 67
        73259 => X"69",  -- 105
        73260 => X"7D",  -- 125
        73261 => X"74",  -- 116
        73262 => X"5B",  -- 91
        73263 => X"60",  -- 96
        73264 => X"5A",  -- 90
        73265 => X"61",  -- 97
        73266 => X"66",  -- 102
        73267 => X"65",  -- 101
        73268 => X"6E",  -- 110
        73269 => X"62",  -- 98
        73270 => X"4D",  -- 77
        73271 => X"5C",  -- 92
        73272 => X"66",  -- 102
        73273 => X"6C",  -- 108
        73274 => X"64",  -- 100
        73275 => X"59",  -- 89
        73276 => X"55",  -- 85
        73277 => X"4D",  -- 77
        73278 => X"47",  -- 71
        73279 => X"4B",  -- 75
        73280 => X"5E",  -- 94
        73281 => X"5B",  -- 91
        73282 => X"5F",  -- 95
        73283 => X"66",  -- 102
        73284 => X"5E",  -- 94
        73285 => X"51",  -- 81
        73286 => X"55",  -- 85
        73287 => X"64",  -- 100
        73288 => X"5C",  -- 92
        73289 => X"5F",  -- 95
        73290 => X"5E",  -- 94
        73291 => X"5A",  -- 90
        73292 => X"5A",  -- 90
        73293 => X"5E",  -- 94
        73294 => X"5C",  -- 92
        73295 => X"57",  -- 87
        73296 => X"50",  -- 80
        73297 => X"54",  -- 84
        73298 => X"59",  -- 89
        73299 => X"5A",  -- 90
        73300 => X"53",  -- 83
        73301 => X"4C",  -- 76
        73302 => X"4E",  -- 78
        73303 => X"55",  -- 85
        73304 => X"4D",  -- 77
        73305 => X"54",  -- 84
        73306 => X"48",  -- 72
        73307 => X"6F",  -- 111
        73308 => X"56",  -- 86
        73309 => X"54",  -- 84
        73310 => X"4E",  -- 78
        73311 => X"45",  -- 69
        73312 => X"50",  -- 80
        73313 => X"4E",  -- 78
        73314 => X"50",  -- 80
        73315 => X"4E",  -- 78
        73316 => X"55",  -- 85
        73317 => X"4F",  -- 79
        73318 => X"49",  -- 73
        73319 => X"69",  -- 105
        73320 => X"52",  -- 82
        73321 => X"48",  -- 72
        73322 => X"42",  -- 66
        73323 => X"56",  -- 86
        73324 => X"5C",  -- 92
        73325 => X"57",  -- 87
        73326 => X"45",  -- 69
        73327 => X"55",  -- 85
        73328 => X"4F",  -- 79
        73329 => X"31",  -- 49
        73330 => X"37",  -- 55
        73331 => X"38",  -- 56
        73332 => X"30",  -- 48
        73333 => X"2D",  -- 45
        73334 => X"3B",  -- 59
        73335 => X"2F",  -- 47
        73336 => X"20",  -- 32
        73337 => X"20",  -- 32
        73338 => X"24",  -- 36
        73339 => X"28",  -- 40
        73340 => X"28",  -- 40
        73341 => X"25",  -- 37
        73342 => X"24",  -- 36
        73343 => X"27",  -- 39
        73344 => X"30",  -- 48
        73345 => X"30",  -- 48
        73346 => X"39",  -- 57
        73347 => X"43",  -- 67
        73348 => X"3E",  -- 62
        73349 => X"2C",  -- 44
        73350 => X"1F",  -- 31
        73351 => X"1D",  -- 29
        73352 => X"21",  -- 33
        73353 => X"39",  -- 57
        73354 => X"49",  -- 73
        73355 => X"42",  -- 66
        73356 => X"2E",  -- 46
        73357 => X"22",  -- 34
        73358 => X"20",  -- 32
        73359 => X"21",  -- 33
        73360 => X"19",  -- 25
        73361 => X"1F",  -- 31
        73362 => X"2E",  -- 46
        73363 => X"37",  -- 55
        73364 => X"37",  -- 55
        73365 => X"37",  -- 55
        73366 => X"33",  -- 51
        73367 => X"26",  -- 38
        73368 => X"1F",  -- 31
        73369 => X"24",  -- 36
        73370 => X"26",  -- 38
        73371 => X"23",  -- 35
        73372 => X"20",  -- 32
        73373 => X"21",  -- 33
        73374 => X"21",  -- 33
        73375 => X"1F",  -- 31
        73376 => X"1D",  -- 29
        73377 => X"1C",  -- 28
        73378 => X"1D",  -- 29
        73379 => X"1D",  -- 29
        73380 => X"1A",  -- 26
        73381 => X"19",  -- 25
        73382 => X"1F",  -- 31
        73383 => X"27",  -- 39
        73384 => X"2D",  -- 45
        73385 => X"28",  -- 40
        73386 => X"25",  -- 37
        73387 => X"24",  -- 36
        73388 => X"1E",  -- 30
        73389 => X"16",  -- 22
        73390 => X"16",  -- 22
        73391 => X"1D",  -- 29
        73392 => X"1B",  -- 27
        73393 => X"1E",  -- 30
        73394 => X"2B",  -- 43
        73395 => X"33",  -- 51
        73396 => X"31",  -- 49
        73397 => X"33",  -- 51
        73398 => X"36",  -- 54
        73399 => X"31",  -- 49
        73400 => X"34",  -- 52
        73401 => X"32",  -- 50
        73402 => X"2E",  -- 46
        73403 => X"2A",  -- 42
        73404 => X"2B",  -- 43
        73405 => X"2E",  -- 46
        73406 => X"2C",  -- 44
        73407 => X"28",  -- 40
        73408 => X"2E",  -- 46
        73409 => X"31",  -- 49
        73410 => X"30",  -- 48
        73411 => X"2A",  -- 42
        73412 => X"28",  -- 40
        73413 => X"2C",  -- 44
        73414 => X"33",  -- 51
        73415 => X"36",  -- 54
        73416 => X"2A",  -- 42
        73417 => X"2E",  -- 46
        73418 => X"33",  -- 51
        73419 => X"35",  -- 53
        73420 => X"34",  -- 52
        73421 => X"34",  -- 52
        73422 => X"34",  -- 52
        73423 => X"35",  -- 53
        73424 => X"33",  -- 51
        73425 => X"2D",  -- 45
        73426 => X"35",  -- 53
        73427 => X"26",  -- 38
        73428 => X"27",  -- 39
        73429 => X"3B",  -- 59
        73430 => X"37",  -- 55
        73431 => X"3E",  -- 62
        73432 => X"41",  -- 65
        73433 => X"4F",  -- 79
        73434 => X"58",  -- 88
        73435 => X"5A",  -- 90
        73436 => X"62",  -- 98
        73437 => X"73",  -- 115
        73438 => X"79",  -- 121
        73439 => X"73",  -- 115
        73440 => X"75",  -- 117
        73441 => X"75",  -- 117
        73442 => X"6A",  -- 106
        73443 => X"6E",  -- 110
        73444 => X"6C",  -- 108
        73445 => X"63",  -- 99
        73446 => X"68",  -- 104
        73447 => X"64",  -- 100
        73448 => X"5C",  -- 92
        73449 => X"5B",  -- 91
        73450 => X"5A",  -- 90
        73451 => X"58",  -- 88
        73452 => X"53",  -- 83
        73453 => X"50",  -- 80
        73454 => X"54",  -- 84
        73455 => X"5A",  -- 90
        73456 => X"6A",  -- 106
        73457 => X"73",  -- 115
        73458 => X"7F",  -- 127
        73459 => X"89",  -- 137
        73460 => X"8E",  -- 142
        73461 => X"87",  -- 135
        73462 => X"6E",  -- 110
        73463 => X"56",  -- 86
        73464 => X"34",  -- 52
        73465 => X"3B",  -- 59
        73466 => X"54",  -- 84
        73467 => X"5E",  -- 94
        73468 => X"4F",  -- 79
        73469 => X"4B",  -- 75
        73470 => X"53",  -- 83
        73471 => X"55",  -- 85
        73472 => X"44",  -- 68
        73473 => X"44",  -- 68
        73474 => X"52",  -- 82
        73475 => X"59",  -- 89
        73476 => X"52",  -- 82
        73477 => X"50",  -- 80
        73478 => X"54",  -- 84
        73479 => X"51",  -- 81
        73480 => X"5E",  -- 94
        73481 => X"5E",  -- 94
        73482 => X"5E",  -- 94
        73483 => X"61",  -- 97
        73484 => X"65",  -- 101
        73485 => X"5E",  -- 94
        73486 => X"59",  -- 89
        73487 => X"63",  -- 99
        73488 => X"68",  -- 104
        73489 => X"6E",  -- 110
        73490 => X"73",  -- 115
        73491 => X"6B",  -- 107
        73492 => X"5F",  -- 95
        73493 => X"58",  -- 88
        73494 => X"5F",  -- 95
        73495 => X"68",  -- 104
        73496 => X"42",  -- 66
        73497 => X"38",  -- 56
        73498 => X"36",  -- 54
        73499 => X"47",  -- 71
        73500 => X"3C",  -- 60
        73501 => X"4C",  -- 76
        73502 => X"35",  -- 53
        73503 => X"32",  -- 50
        73504 => X"51",  -- 81
        73505 => X"52",  -- 82
        73506 => X"51",  -- 81
        73507 => X"4F",  -- 79
        73508 => X"4D",  -- 77
        73509 => X"4A",  -- 74
        73510 => X"47",  -- 71
        73511 => X"42",  -- 66
        73512 => X"40",  -- 64
        73513 => X"48",  -- 72
        73514 => X"4E",  -- 78
        73515 => X"4E",  -- 78
        73516 => X"54",  -- 84
        73517 => X"56",  -- 86
        73518 => X"4F",  -- 79
        73519 => X"41",  -- 65
        73520 => X"3A",  -- 58
        73521 => X"50",  -- 80
        73522 => X"5A",  -- 90
        73523 => X"55",  -- 85
        73524 => X"53",  -- 83
        73525 => X"57",  -- 87
        73526 => X"5C",  -- 92
        73527 => X"60",  -- 96
        73528 => X"5E",  -- 94
        73529 => X"6A",  -- 106
        73530 => X"63",  -- 99
        73531 => X"58",  -- 88
        73532 => X"57",  -- 87
        73533 => X"65",  -- 101
        73534 => X"5C",  -- 92
        73535 => X"68",  -- 104
        73536 => X"6E",  -- 110
        73537 => X"64",  -- 100
        73538 => X"63",  -- 99
        73539 => X"72",  -- 114
        73540 => X"7B",  -- 123
        73541 => X"74",  -- 116
        73542 => X"71",  -- 113
        73543 => X"77",  -- 119
        73544 => X"59",  -- 89
        73545 => X"5D",  -- 93
        73546 => X"48",  -- 72
        73547 => X"43",  -- 67
        73548 => X"5C",  -- 92
        73549 => X"72",  -- 114
        73550 => X"6B",  -- 107
        73551 => X"63",  -- 99
        73552 => X"6A",  -- 106
        73553 => X"60",  -- 96
        73554 => X"60",  -- 96
        73555 => X"58",  -- 88
        73556 => X"66",  -- 102
        73557 => X"8D",  -- 141
        73558 => X"99",  -- 153
        73559 => X"9B",  -- 155
        73560 => X"9A",  -- 154
        73561 => X"A6",  -- 166
        73562 => X"9F",  -- 159
        73563 => X"A3",  -- 163
        73564 => X"A9",  -- 169
        73565 => X"5A",  -- 90
        73566 => X"5A",  -- 90
        73567 => X"4B",  -- 75
        73568 => X"5C",  -- 92
        73569 => X"5C",  -- 92
        73570 => X"53",  -- 83
        73571 => X"63",  -- 99
        73572 => X"44",  -- 68
        73573 => X"43",  -- 67
        73574 => X"5E",  -- 94
        73575 => X"5D",  -- 93
        73576 => X"43",  -- 67
        73577 => X"25",  -- 37
        73578 => X"34",  -- 52
        73579 => X"48",  -- 72
        73580 => X"63",  -- 99
        73581 => X"74",  -- 116
        73582 => X"54",  -- 84
        73583 => X"42",  -- 66
        73584 => X"6D",  -- 109
        73585 => X"4C",  -- 76
        73586 => X"63",  -- 99
        73587 => X"75",  -- 117
        73588 => X"6F",  -- 111
        73589 => X"72",  -- 114
        73590 => X"60",  -- 96
        73591 => X"45",  -- 69
        73592 => X"6A",  -- 106
        73593 => X"76",  -- 118
        73594 => X"72",  -- 114
        73595 => X"66",  -- 102
        73596 => X"60",  -- 96
        73597 => X"59",  -- 89
        73598 => X"52",  -- 82
        73599 => X"52",  -- 82
        73600 => X"5B",  -- 91
        73601 => X"59",  -- 89
        73602 => X"5D",  -- 93
        73603 => X"63",  -- 99
        73604 => X"5C",  -- 92
        73605 => X"50",  -- 80
        73606 => X"56",  -- 86
        73607 => X"66",  -- 102
        73608 => X"58",  -- 88
        73609 => X"5B",  -- 91
        73610 => X"5D",  -- 93
        73611 => X"5E",  -- 94
        73612 => X"5E",  -- 94
        73613 => X"5D",  -- 93
        73614 => X"5A",  -- 90
        73615 => X"57",  -- 87
        73616 => X"52",  -- 82
        73617 => X"5C",  -- 92
        73618 => X"64",  -- 100
        73619 => X"5F",  -- 95
        73620 => X"57",  -- 87
        73621 => X"54",  -- 84
        73622 => X"56",  -- 86
        73623 => X"57",  -- 87
        73624 => X"46",  -- 70
        73625 => X"46",  -- 70
        73626 => X"46",  -- 70
        73627 => X"73",  -- 115
        73628 => X"41",  -- 65
        73629 => X"57",  -- 87
        73630 => X"55",  -- 85
        73631 => X"52",  -- 82
        73632 => X"4D",  -- 77
        73633 => X"45",  -- 69
        73634 => X"43",  -- 67
        73635 => X"45",  -- 69
        73636 => X"51",  -- 81
        73637 => X"4D",  -- 77
        73638 => X"51",  -- 81
        73639 => X"81",  -- 129
        73640 => X"51",  -- 81
        73641 => X"46",  -- 70
        73642 => X"3E",  -- 62
        73643 => X"32",  -- 50
        73644 => X"44",  -- 68
        73645 => X"41",  -- 65
        73646 => X"38",  -- 56
        73647 => X"41",  -- 65
        73648 => X"4F",  -- 79
        73649 => X"2A",  -- 42
        73650 => X"38",  -- 56
        73651 => X"42",  -- 66
        73652 => X"3F",  -- 63
        73653 => X"34",  -- 52
        73654 => X"40",  -- 64
        73655 => X"30",  -- 48
        73656 => X"20",  -- 32
        73657 => X"1F",  -- 31
        73658 => X"21",  -- 33
        73659 => X"26",  -- 38
        73660 => X"29",  -- 41
        73661 => X"2A",  -- 42
        73662 => X"2D",  -- 45
        73663 => X"31",  -- 49
        73664 => X"3B",  -- 59
        73665 => X"34",  -- 52
        73666 => X"39",  -- 57
        73667 => X"45",  -- 69
        73668 => X"3F",  -- 63
        73669 => X"27",  -- 39
        73670 => X"1C",  -- 28
        73671 => X"20",  -- 32
        73672 => X"25",  -- 37
        73673 => X"3A",  -- 58
        73674 => X"49",  -- 73
        73675 => X"43",  -- 67
        73676 => X"33",  -- 51
        73677 => X"28",  -- 40
        73678 => X"20",  -- 32
        73679 => X"1B",  -- 27
        73680 => X"1B",  -- 27
        73681 => X"21",  -- 33
        73682 => X"2E",  -- 46
        73683 => X"35",  -- 53
        73684 => X"35",  -- 53
        73685 => X"39",  -- 57
        73686 => X"3A",  -- 58
        73687 => X"30",  -- 48
        73688 => X"1F",  -- 31
        73689 => X"21",  -- 33
        73690 => X"20",  -- 32
        73691 => X"1E",  -- 30
        73692 => X"1E",  -- 30
        73693 => X"20",  -- 32
        73694 => X"1F",  -- 31
        73695 => X"1C",  -- 28
        73696 => X"1F",  -- 31
        73697 => X"1E",  -- 30
        73698 => X"1F",  -- 31
        73699 => X"1F",  -- 31
        73700 => X"1D",  -- 29
        73701 => X"1D",  -- 29
        73702 => X"24",  -- 36
        73703 => X"2D",  -- 45
        73704 => X"35",  -- 53
        73705 => X"30",  -- 48
        73706 => X"2D",  -- 45
        73707 => X"2B",  -- 43
        73708 => X"23",  -- 35
        73709 => X"18",  -- 24
        73710 => X"17",  -- 23
        73711 => X"1E",  -- 30
        73712 => X"1C",  -- 28
        73713 => X"1A",  -- 26
        73714 => X"28",  -- 40
        73715 => X"37",  -- 55
        73716 => X"35",  -- 53
        73717 => X"30",  -- 48
        73718 => X"32",  -- 50
        73719 => X"31",  -- 49
        73720 => X"33",  -- 51
        73721 => X"31",  -- 49
        73722 => X"2C",  -- 44
        73723 => X"27",  -- 39
        73724 => X"28",  -- 40
        73725 => X"2E",  -- 46
        73726 => X"2F",  -- 47
        73727 => X"2D",  -- 45
        73728 => X"2D",  -- 45
        73729 => X"30",  -- 48
        73730 => X"30",  -- 48
        73731 => X"2B",  -- 43
        73732 => X"29",  -- 41
        73733 => X"2C",  -- 44
        73734 => X"2E",  -- 46
        73735 => X"2C",  -- 44
        73736 => X"26",  -- 38
        73737 => X"2A",  -- 42
        73738 => X"33",  -- 51
        73739 => X"39",  -- 57
        73740 => X"3D",  -- 61
        73741 => X"3C",  -- 60
        73742 => X"3A",  -- 58
        73743 => X"38",  -- 56
        73744 => X"38",  -- 56
        73745 => X"33",  -- 51
        73746 => X"35",  -- 53
        73747 => X"2E",  -- 46
        73748 => X"33",  -- 51
        73749 => X"4B",  -- 75
        73750 => X"55",  -- 85
        73751 => X"56",  -- 86
        73752 => X"4F",  -- 79
        73753 => X"62",  -- 98
        73754 => X"6D",  -- 109
        73755 => X"6B",  -- 107
        73756 => X"69",  -- 105
        73757 => X"6A",  -- 106
        73758 => X"6B",  -- 107
        73759 => X"70",  -- 112
        73760 => X"68",  -- 104
        73761 => X"61",  -- 97
        73762 => X"55",  -- 85
        73763 => X"5B",  -- 91
        73764 => X"57",  -- 87
        73765 => X"47",  -- 71
        73766 => X"4C",  -- 76
        73767 => X"4E",  -- 78
        73768 => X"45",  -- 69
        73769 => X"41",  -- 65
        73770 => X"40",  -- 64
        73771 => X"40",  -- 64
        73772 => X"3F",  -- 63
        73773 => X"3B",  -- 59
        73774 => X"3A",  -- 58
        73775 => X"3D",  -- 61
        73776 => X"4D",  -- 77
        73777 => X"54",  -- 84
        73778 => X"61",  -- 97
        73779 => X"74",  -- 116
        73780 => X"83",  -- 131
        73781 => X"83",  -- 131
        73782 => X"77",  -- 119
        73783 => X"6A",  -- 106
        73784 => X"4C",  -- 76
        73785 => X"43",  -- 67
        73786 => X"4B",  -- 75
        73787 => X"60",  -- 96
        73788 => X"61",  -- 97
        73789 => X"52",  -- 82
        73790 => X"4C",  -- 76
        73791 => X"51",  -- 81
        73792 => X"41",  -- 65
        73793 => X"39",  -- 57
        73794 => X"45",  -- 69
        73795 => X"51",  -- 81
        73796 => X"4C",  -- 76
        73797 => X"4E",  -- 78
        73798 => X"53",  -- 83
        73799 => X"4F",  -- 79
        73800 => X"57",  -- 87
        73801 => X"5E",  -- 94
        73802 => X"61",  -- 97
        73803 => X"63",  -- 99
        73804 => X"67",  -- 103
        73805 => X"62",  -- 98
        73806 => X"5C",  -- 92
        73807 => X"5F",  -- 95
        73808 => X"5F",  -- 95
        73809 => X"66",  -- 102
        73810 => X"65",  -- 101
        73811 => X"5D",  -- 93
        73812 => X"58",  -- 88
        73813 => X"5E",  -- 94
        73814 => X"63",  -- 99
        73815 => X"64",  -- 100
        73816 => X"58",  -- 88
        73817 => X"49",  -- 73
        73818 => X"49",  -- 73
        73819 => X"54",  -- 84
        73820 => X"45",  -- 69
        73821 => X"52",  -- 82
        73822 => X"43",  -- 67
        73823 => X"40",  -- 64
        73824 => X"55",  -- 85
        73825 => X"54",  -- 84
        73826 => X"51",  -- 81
        73827 => X"4A",  -- 74
        73828 => X"48",  -- 72
        73829 => X"49",  -- 73
        73830 => X"46",  -- 70
        73831 => X"41",  -- 65
        73832 => X"44",  -- 68
        73833 => X"48",  -- 72
        73834 => X"4E",  -- 78
        73835 => X"4F",  -- 79
        73836 => X"4E",  -- 78
        73837 => X"4D",  -- 77
        73838 => X"49",  -- 73
        73839 => X"43",  -- 67
        73840 => X"45",  -- 69
        73841 => X"4C",  -- 76
        73842 => X"5D",  -- 93
        73843 => X"62",  -- 98
        73844 => X"54",  -- 84
        73845 => X"46",  -- 70
        73846 => X"43",  -- 67
        73847 => X"44",  -- 68
        73848 => X"41",  -- 65
        73849 => X"72",  -- 114
        73850 => X"6E",  -- 110
        73851 => X"61",  -- 97
        73852 => X"58",  -- 88
        73853 => X"69",  -- 105
        73854 => X"66",  -- 102
        73855 => X"5E",  -- 94
        73856 => X"5D",  -- 93
        73857 => X"61",  -- 97
        73858 => X"64",  -- 100
        73859 => X"6B",  -- 107
        73860 => X"70",  -- 112
        73861 => X"6F",  -- 111
        73862 => X"6D",  -- 109
        73863 => X"72",  -- 114
        73864 => X"4D",  -- 77
        73865 => X"56",  -- 86
        73866 => X"5D",  -- 93
        73867 => X"59",  -- 89
        73868 => X"61",  -- 97
        73869 => X"72",  -- 114
        73870 => X"6A",  -- 106
        73871 => X"4B",  -- 75
        73872 => X"5D",  -- 93
        73873 => X"57",  -- 87
        73874 => X"4B",  -- 75
        73875 => X"57",  -- 87
        73876 => X"8C",  -- 140
        73877 => X"A5",  -- 165
        73878 => X"98",  -- 152
        73879 => X"AA",  -- 170
        73880 => X"9C",  -- 156
        73881 => X"9A",  -- 154
        73882 => X"93",  -- 147
        73883 => X"8C",  -- 140
        73884 => X"84",  -- 132
        73885 => X"60",  -- 96
        73886 => X"72",  -- 114
        73887 => X"6C",  -- 108
        73888 => X"68",  -- 104
        73889 => X"64",  -- 100
        73890 => X"4F",  -- 79
        73891 => X"67",  -- 103
        73892 => X"44",  -- 68
        73893 => X"26",  -- 38
        73894 => X"37",  -- 55
        73895 => X"45",  -- 69
        73896 => X"43",  -- 67
        73897 => X"26",  -- 38
        73898 => X"2F",  -- 47
        73899 => X"2E",  -- 46
        73900 => X"46",  -- 70
        73901 => X"6E",  -- 110
        73902 => X"59",  -- 89
        73903 => X"43",  -- 67
        73904 => X"50",  -- 80
        73905 => X"48",  -- 72
        73906 => X"61",  -- 97
        73907 => X"7B",  -- 123
        73908 => X"66",  -- 102
        73909 => X"5C",  -- 92
        73910 => X"6A",  -- 106
        73911 => X"53",  -- 83
        73912 => X"62",  -- 98
        73913 => X"74",  -- 116
        73914 => X"77",  -- 119
        73915 => X"6E",  -- 110
        73916 => X"69",  -- 105
        73917 => X"66",  -- 102
        73918 => X"63",  -- 99
        73919 => X"65",  -- 101
        73920 => X"59",  -- 89
        73921 => X"5A",  -- 90
        73922 => X"5F",  -- 95
        73923 => X"63",  -- 99
        73924 => X"5E",  -- 94
        73925 => X"55",  -- 85
        73926 => X"57",  -- 87
        73927 => X"61",  -- 97
        73928 => X"5B",  -- 91
        73929 => X"5D",  -- 93
        73930 => X"62",  -- 98
        73931 => X"64",  -- 100
        73932 => X"61",  -- 97
        73933 => X"5B",  -- 91
        73934 => X"59",  -- 89
        73935 => X"59",  -- 89
        73936 => X"56",  -- 86
        73937 => X"64",  -- 100
        73938 => X"6D",  -- 109
        73939 => X"65",  -- 101
        73940 => X"5B",  -- 91
        73941 => X"5A",  -- 90
        73942 => X"5A",  -- 90
        73943 => X"58",  -- 88
        73944 => X"5E",  -- 94
        73945 => X"4B",  -- 75
        73946 => X"56",  -- 86
        73947 => X"88",  -- 136
        73948 => X"42",  -- 66
        73949 => X"4A",  -- 74
        73950 => X"44",  -- 68
        73951 => X"4A",  -- 74
        73952 => X"48",  -- 72
        73953 => X"42",  -- 66
        73954 => X"41",  -- 65
        73955 => X"41",  -- 65
        73956 => X"46",  -- 70
        73957 => X"3C",  -- 60
        73958 => X"4B",  -- 75
        73959 => X"8B",  -- 139
        73960 => X"4B",  -- 75
        73961 => X"3F",  -- 63
        73962 => X"46",  -- 70
        73963 => X"29",  -- 41
        73964 => X"3F",  -- 63
        73965 => X"37",  -- 55
        73966 => X"1E",  -- 30
        73967 => X"1B",  -- 27
        73968 => X"53",  -- 83
        73969 => X"28",  -- 40
        73970 => X"38",  -- 56
        73971 => X"49",  -- 73
        73972 => X"4C",  -- 76
        73973 => X"3F",  -- 63
        73974 => X"4C",  -- 76
        73975 => X"3A",  -- 58
        73976 => X"20",  -- 32
        73977 => X"1D",  -- 29
        73978 => X"1F",  -- 31
        73979 => X"25",  -- 37
        73980 => X"2B",  -- 43
        73981 => X"30",  -- 48
        73982 => X"38",  -- 56
        73983 => X"3F",  -- 63
        73984 => X"44",  -- 68
        73985 => X"43",  -- 67
        73986 => X"44",  -- 68
        73987 => X"44",  -- 68
        73988 => X"3E",  -- 62
        73989 => X"33",  -- 51
        73990 => X"28",  -- 40
        73991 => X"24",  -- 36
        73992 => X"2B",  -- 43
        73993 => X"3D",  -- 61
        73994 => X"48",  -- 72
        73995 => X"42",  -- 66
        73996 => X"36",  -- 54
        73997 => X"2D",  -- 45
        73998 => X"22",  -- 34
        73999 => X"18",  -- 24
        74000 => X"1E",  -- 30
        74001 => X"26",  -- 38
        74002 => X"34",  -- 52
        74003 => X"39",  -- 57
        74004 => X"36",  -- 54
        74005 => X"39",  -- 57
        74006 => X"3B",  -- 59
        74007 => X"33",  -- 51
        74008 => X"1E",  -- 30
        74009 => X"1F",  -- 31
        74010 => X"1D",  -- 29
        74011 => X"1C",  -- 28
        74012 => X"1F",  -- 31
        74013 => X"23",  -- 35
        74014 => X"22",  -- 34
        74015 => X"1E",  -- 30
        74016 => X"1E",  -- 30
        74017 => X"1D",  -- 29
        74018 => X"1E",  -- 30
        74019 => X"1E",  -- 30
        74020 => X"1B",  -- 27
        74021 => X"1B",  -- 27
        74022 => X"22",  -- 34
        74023 => X"2B",  -- 43
        74024 => X"36",  -- 54
        74025 => X"33",  -- 51
        74026 => X"32",  -- 50
        74027 => X"2F",  -- 47
        74028 => X"25",  -- 37
        74029 => X"18",  -- 24
        74030 => X"16",  -- 22
        74031 => X"1C",  -- 28
        74032 => X"19",  -- 25
        74033 => X"14",  -- 20
        74034 => X"24",  -- 36
        74035 => X"38",  -- 56
        74036 => X"36",  -- 54
        74037 => X"2D",  -- 45
        74038 => X"2D",  -- 45
        74039 => X"2E",  -- 46
        74040 => X"33",  -- 51
        74041 => X"31",  -- 49
        74042 => X"2B",  -- 43
        74043 => X"25",  -- 37
        74044 => X"25",  -- 37
        74045 => X"2B",  -- 43
        74046 => X"2D",  -- 45
        74047 => X"2A",  -- 42
        74048 => X"24",  -- 36
        74049 => X"2A",  -- 42
        74050 => X"2E",  -- 46
        74051 => X"2E",  -- 46
        74052 => X"2F",  -- 47
        74053 => X"33",  -- 51
        74054 => X"32",  -- 50
        74055 => X"2E",  -- 46
        74056 => X"30",  -- 48
        74057 => X"2F",  -- 47
        74058 => X"2E",  -- 46
        74059 => X"2D",  -- 45
        74060 => X"32",  -- 50
        74061 => X"36",  -- 54
        74062 => X"37",  -- 55
        74063 => X"38",  -- 56
        74064 => X"45",  -- 69
        74065 => X"46",  -- 70
        74066 => X"4A",  -- 74
        74067 => X"4B",  -- 75
        74068 => X"4F",  -- 79
        74069 => X"5B",  -- 91
        74070 => X"64",  -- 100
        74071 => X"5C",  -- 92
        74072 => X"60",  -- 96
        74073 => X"61",  -- 97
        74074 => X"60",  -- 96
        74075 => X"67",  -- 103
        74076 => X"6E",  -- 110
        74077 => X"63",  -- 99
        74078 => X"54",  -- 84
        74079 => X"52",  -- 82
        74080 => X"4B",  -- 75
        74081 => X"44",  -- 68
        74082 => X"3C",  -- 60
        74083 => X"49",  -- 73
        74084 => X"46",  -- 70
        74085 => X"35",  -- 53
        74086 => X"3D",  -- 61
        74087 => X"47",  -- 71
        74088 => X"43",  -- 67
        74089 => X"3C",  -- 60
        74090 => X"38",  -- 56
        74091 => X"3C",  -- 60
        74092 => X"3E",  -- 62
        74093 => X"3B",  -- 59
        74094 => X"37",  -- 55
        74095 => X"36",  -- 54
        74096 => X"3A",  -- 58
        74097 => X"3C",  -- 60
        74098 => X"4A",  -- 74
        74099 => X"60",  -- 96
        74100 => X"73",  -- 115
        74101 => X"7A",  -- 122
        74102 => X"7A",  -- 122
        74103 => X"77",  -- 119
        74104 => X"6A",  -- 106
        74105 => X"50",  -- 80
        74106 => X"45",  -- 69
        74107 => X"5D",  -- 93
        74108 => X"6B",  -- 107
        74109 => X"53",  -- 83
        74110 => X"40",  -- 64
        74111 => X"47",  -- 71
        74112 => X"40",  -- 64
        74113 => X"33",  -- 51
        74114 => X"3A",  -- 58
        74115 => X"48",  -- 72
        74116 => X"47",  -- 71
        74117 => X"4C",  -- 76
        74118 => X"54",  -- 84
        74119 => X"4C",  -- 76
        74120 => X"4F",  -- 79
        74121 => X"5E",  -- 94
        74122 => X"62",  -- 98
        74123 => X"65",  -- 101
        74124 => X"6B",  -- 107
        74125 => X"69",  -- 105
        74126 => X"63",  -- 99
        74127 => X"62",  -- 98
        74128 => X"6A",  -- 106
        74129 => X"68",  -- 104
        74130 => X"5E",  -- 94
        74131 => X"56",  -- 86
        74132 => X"5E",  -- 94
        74133 => X"68",  -- 104
        74134 => X"5F",  -- 95
        74135 => X"4C",  -- 76
        74136 => X"57",  -- 87
        74137 => X"3F",  -- 63
        74138 => X"52",  -- 82
        74139 => X"47",  -- 71
        74140 => X"4D",  -- 77
        74141 => X"49",  -- 73
        74142 => X"52",  -- 82
        74143 => X"4C",  -- 76
        74144 => X"42",  -- 66
        74145 => X"4B",  -- 75
        74146 => X"51",  -- 81
        74147 => X"4B",  -- 75
        74148 => X"44",  -- 68
        74149 => X"45",  -- 69
        74150 => X"44",  -- 68
        74151 => X"43",  -- 67
        74152 => X"4C",  -- 76
        74153 => X"4A",  -- 74
        74154 => X"4A",  -- 74
        74155 => X"4D",  -- 77
        74156 => X"48",  -- 72
        74157 => X"41",  -- 65
        74158 => X"45",  -- 69
        74159 => X"4D",  -- 77
        74160 => X"53",  -- 83
        74161 => X"3D",  -- 61
        74162 => X"43",  -- 67
        74163 => X"55",  -- 85
        74164 => X"4F",  -- 79
        74165 => X"48",  -- 72
        74166 => X"50",  -- 80
        74167 => X"57",  -- 87
        74168 => X"50",  -- 80
        74169 => X"59",  -- 89
        74170 => X"5D",  -- 93
        74171 => X"7A",  -- 122
        74172 => X"63",  -- 99
        74173 => X"6D",  -- 109
        74174 => X"73",  -- 115
        74175 => X"4F",  -- 79
        74176 => X"2D",  -- 45
        74177 => X"59",  -- 89
        74178 => X"6F",  -- 111
        74179 => X"67",  -- 103
        74180 => X"6A",  -- 106
        74181 => X"73",  -- 115
        74182 => X"6B",  -- 107
        74183 => X"5C",  -- 92
        74184 => X"59",  -- 89
        74185 => X"3E",  -- 62
        74186 => X"5A",  -- 90
        74187 => X"7B",  -- 123
        74188 => X"6F",  -- 111
        74189 => X"64",  -- 100
        74190 => X"69",  -- 105
        74191 => X"5A",  -- 90
        74192 => X"61",  -- 97
        74193 => X"31",  -- 49
        74194 => X"41",  -- 65
        74195 => X"75",  -- 117
        74196 => X"8E",  -- 142
        74197 => X"94",  -- 148
        74198 => X"94",  -- 148
        74199 => X"A4",  -- 164
        74200 => X"9E",  -- 158
        74201 => X"94",  -- 148
        74202 => X"A4",  -- 164
        74203 => X"9F",  -- 159
        74204 => X"79",  -- 121
        74205 => X"6F",  -- 111
        74206 => X"75",  -- 117
        74207 => X"69",  -- 105
        74208 => X"5E",  -- 94
        74209 => X"73",  -- 115
        74210 => X"58",  -- 88
        74211 => X"57",  -- 87
        74212 => X"36",  -- 54
        74213 => X"22",  -- 34
        74214 => X"2C",  -- 44
        74215 => X"26",  -- 38
        74216 => X"2F",  -- 47
        74217 => X"1D",  -- 29
        74218 => X"37",  -- 55
        74219 => X"37",  -- 55
        74220 => X"42",  -- 66
        74221 => X"63",  -- 99
        74222 => X"53",  -- 83
        74223 => X"46",  -- 70
        74224 => X"47",  -- 71
        74225 => X"57",  -- 87
        74226 => X"44",  -- 68
        74227 => X"68",  -- 104
        74228 => X"7D",  -- 125
        74229 => X"68",  -- 104
        74230 => X"71",  -- 113
        74231 => X"5C",  -- 92
        74232 => X"62",  -- 98
        74233 => X"76",  -- 118
        74234 => X"79",  -- 121
        74235 => X"6E",  -- 110
        74236 => X"69",  -- 105
        74237 => X"69",  -- 105
        74238 => X"6A",  -- 106
        74239 => X"6D",  -- 109
        74240 => X"51",  -- 81
        74241 => X"56",  -- 86
        74242 => X"63",  -- 99
        74243 => X"69",  -- 105
        74244 => X"62",  -- 98
        74245 => X"60",  -- 96
        74246 => X"62",  -- 98
        74247 => X"5E",  -- 94
        74248 => X"64",  -- 100
        74249 => X"5B",  -- 91
        74250 => X"5B",  -- 91
        74251 => X"65",  -- 101
        74252 => X"66",  -- 102
        74253 => X"5B",  -- 91
        74254 => X"56",  -- 86
        74255 => X"59",  -- 89
        74256 => X"61",  -- 97
        74257 => X"65",  -- 101
        74258 => X"61",  -- 97
        74259 => X"5E",  -- 94
        74260 => X"5E",  -- 94
        74261 => X"55",  -- 85
        74262 => X"49",  -- 73
        74263 => X"48",  -- 72
        74264 => X"34",  -- 52
        74265 => X"47",  -- 71
        74266 => X"5E",  -- 94
        74267 => X"72",  -- 114
        74268 => X"5C",  -- 92
        74269 => X"44",  -- 68
        74270 => X"48",  -- 72
        74271 => X"4C",  -- 76
        74272 => X"50",  -- 80
        74273 => X"4D",  -- 77
        74274 => X"4D",  -- 77
        74275 => X"4A",  -- 74
        74276 => X"3B",  -- 59
        74277 => X"36",  -- 54
        74278 => X"4F",  -- 79
        74279 => X"70",  -- 112
        74280 => X"43",  -- 67
        74281 => X"39",  -- 57
        74282 => X"35",  -- 53
        74283 => X"26",  -- 38
        74284 => X"4A",  -- 74
        74285 => X"26",  -- 38
        74286 => X"1C",  -- 28
        74287 => X"1E",  -- 30
        74288 => X"2C",  -- 44
        74289 => X"55",  -- 85
        74290 => X"41",  -- 65
        74291 => X"47",  -- 71
        74292 => X"46",  -- 70
        74293 => X"44",  -- 68
        74294 => X"38",  -- 56
        74295 => X"33",  -- 51
        74296 => X"1B",  -- 27
        74297 => X"29",  -- 41
        74298 => X"2C",  -- 44
        74299 => X"29",  -- 41
        74300 => X"28",  -- 40
        74301 => X"27",  -- 39
        74302 => X"2D",  -- 45
        74303 => X"3B",  -- 59
        74304 => X"43",  -- 67
        74305 => X"47",  -- 71
        74306 => X"42",  -- 66
        74307 => X"3E",  -- 62
        74308 => X"3E",  -- 62
        74309 => X"33",  -- 51
        74310 => X"25",  -- 37
        74311 => X"21",  -- 33
        74312 => X"2B",  -- 43
        74313 => X"4C",  -- 76
        74314 => X"4C",  -- 76
        74315 => X"3B",  -- 59
        74316 => X"3C",  -- 60
        74317 => X"30",  -- 48
        74318 => X"1C",  -- 28
        74319 => X"1B",  -- 27
        74320 => X"23",  -- 35
        74321 => X"2F",  -- 47
        74322 => X"38",  -- 56
        74323 => X"37",  -- 55
        74324 => X"33",  -- 51
        74325 => X"32",  -- 50
        74326 => X"33",  -- 51
        74327 => X"33",  -- 51
        74328 => X"1C",  -- 28
        74329 => X"23",  -- 35
        74330 => X"21",  -- 33
        74331 => X"1E",  -- 30
        74332 => X"22",  -- 34
        74333 => X"21",  -- 33
        74334 => X"1D",  -- 29
        74335 => X"1F",  -- 31
        74336 => X"24",  -- 36
        74337 => X"20",  -- 32
        74338 => X"21",  -- 33
        74339 => X"19",  -- 25
        74340 => X"19",  -- 25
        74341 => X"1C",  -- 28
        74342 => X"22",  -- 34
        74343 => X"3D",  -- 61
        74344 => X"39",  -- 57
        74345 => X"3E",  -- 62
        74346 => X"34",  -- 52
        74347 => X"24",  -- 36
        74348 => X"1C",  -- 28
        74349 => X"17",  -- 23
        74350 => X"14",  -- 20
        74351 => X"19",  -- 25
        74352 => X"18",  -- 24
        74353 => X"1F",  -- 31
        74354 => X"25",  -- 37
        74355 => X"2E",  -- 46
        74356 => X"35",  -- 53
        74357 => X"2F",  -- 47
        74358 => X"29",  -- 41
        74359 => X"2F",  -- 47
        74360 => X"33",  -- 51
        74361 => X"2D",  -- 45
        74362 => X"2B",  -- 43
        74363 => X"2E",  -- 46
        74364 => X"2B",  -- 43
        74365 => X"26",  -- 38
        74366 => X"2A",  -- 42
        74367 => X"35",  -- 53
        74368 => X"30",  -- 48
        74369 => X"2E",  -- 46
        74370 => X"2A",  -- 42
        74371 => X"2C",  -- 44
        74372 => X"2D",  -- 45
        74373 => X"2F",  -- 47
        74374 => X"30",  -- 48
        74375 => X"2E",  -- 46
        74376 => X"1E",  -- 30
        74377 => X"2E",  -- 46
        74378 => X"37",  -- 55
        74379 => X"32",  -- 50
        74380 => X"2F",  -- 47
        74381 => X"39",  -- 57
        74382 => X"43",  -- 67
        74383 => X"47",  -- 71
        74384 => X"52",  -- 82
        74385 => X"51",  -- 81
        74386 => X"5D",  -- 93
        74387 => X"61",  -- 97
        74388 => X"58",  -- 88
        74389 => X"5F",  -- 95
        74390 => X"66",  -- 102
        74391 => X"5A",  -- 90
        74392 => X"56",  -- 86
        74393 => X"65",  -- 101
        74394 => X"60",  -- 96
        74395 => X"57",  -- 87
        74396 => X"56",  -- 86
        74397 => X"46",  -- 70
        74398 => X"2F",  -- 47
        74399 => X"2A",  -- 42
        74400 => X"33",  -- 51
        74401 => X"32",  -- 50
        74402 => X"2D",  -- 45
        74403 => X"29",  -- 41
        74404 => X"35",  -- 53
        74405 => X"42",  -- 66
        74406 => X"3F",  -- 63
        74407 => X"33",  -- 51
        74408 => X"39",  -- 57
        74409 => X"3C",  -- 60
        74410 => X"44",  -- 68
        74411 => X"42",  -- 66
        74412 => X"3F",  -- 63
        74413 => X"46",  -- 70
        74414 => X"49",  -- 73
        74415 => X"3E",  -- 62
        74416 => X"36",  -- 54
        74417 => X"31",  -- 49
        74418 => X"2C",  -- 44
        74419 => X"39",  -- 57
        74420 => X"5A",  -- 90
        74421 => X"6F",  -- 111
        74422 => X"72",  -- 114
        74423 => X"75",  -- 117
        74424 => X"6C",  -- 108
        74425 => X"56",  -- 86
        74426 => X"51",  -- 81
        74427 => X"63",  -- 99
        74428 => X"64",  -- 100
        74429 => X"4E",  -- 78
        74430 => X"44",  -- 68
        74431 => X"4F",  -- 79
        74432 => X"34",  -- 52
        74433 => X"38",  -- 56
        74434 => X"3F",  -- 63
        74435 => X"47",  -- 71
        74436 => X"4C",  -- 76
        74437 => X"4D",  -- 77
        74438 => X"4F",  -- 79
        74439 => X"4F",  -- 79
        74440 => X"4A",  -- 74
        74441 => X"51",  -- 81
        74442 => X"5A",  -- 90
        74443 => X"60",  -- 96
        74444 => X"64",  -- 100
        74445 => X"66",  -- 102
        74446 => X"6A",  -- 106
        74447 => X"6E",  -- 110
        74448 => X"69",  -- 105
        74449 => X"5F",  -- 95
        74450 => X"5C",  -- 92
        74451 => X"5D",  -- 93
        74452 => X"56",  -- 86
        74453 => X"4B",  -- 75
        74454 => X"58",  -- 88
        74455 => X"6D",  -- 109
        74456 => X"64",  -- 100
        74457 => X"40",  -- 64
        74458 => X"45",  -- 69
        74459 => X"45",  -- 69
        74460 => X"41",  -- 65
        74461 => X"4B",  -- 75
        74462 => X"44",  -- 68
        74463 => X"48",  -- 72
        74464 => X"3B",  -- 59
        74465 => X"42",  -- 66
        74466 => X"4A",  -- 74
        74467 => X"4C",  -- 76
        74468 => X"47",  -- 71
        74469 => X"41",  -- 65
        74470 => X"3F",  -- 63
        74471 => X"41",  -- 65
        74472 => X"49",  -- 73
        74473 => X"4A",  -- 74
        74474 => X"4B",  -- 75
        74475 => X"4F",  -- 79
        74476 => X"55",  -- 85
        74477 => X"59",  -- 89
        74478 => X"55",  -- 85
        74479 => X"50",  -- 80
        74480 => X"59",  -- 89
        74481 => X"54",  -- 84
        74482 => X"47",  -- 71
        74483 => X"44",  -- 68
        74484 => X"4C",  -- 76
        74485 => X"4B",  -- 75
        74486 => X"43",  -- 67
        74487 => X"44",  -- 68
        74488 => X"4F",  -- 79
        74489 => X"3F",  -- 63
        74490 => X"56",  -- 86
        74491 => X"63",  -- 99
        74492 => X"79",  -- 121
        74493 => X"6D",  -- 109
        74494 => X"67",  -- 103
        74495 => X"6B",  -- 107
        74496 => X"98",  -- 152
        74497 => X"78",  -- 120
        74498 => X"6E",  -- 110
        74499 => X"6C",  -- 108
        74500 => X"60",  -- 96
        74501 => X"5E",  -- 94
        74502 => X"5B",  -- 91
        74503 => X"4A",  -- 74
        74504 => X"3F",  -- 63
        74505 => X"3F",  -- 63
        74506 => X"5B",  -- 91
        74507 => X"81",  -- 129
        74508 => X"58",  -- 88
        74509 => X"57",  -- 87
        74510 => X"73",  -- 115
        74511 => X"9A",  -- 154
        74512 => X"49",  -- 73
        74513 => X"33",  -- 51
        74514 => X"53",  -- 83
        74515 => X"6C",  -- 108
        74516 => X"99",  -- 153
        74517 => X"8A",  -- 138
        74518 => X"93",  -- 147
        74519 => X"9A",  -- 154
        74520 => X"90",  -- 144
        74521 => X"9E",  -- 158
        74522 => X"8C",  -- 140
        74523 => X"85",  -- 133
        74524 => X"7D",  -- 125
        74525 => X"56",  -- 86
        74526 => X"72",  -- 114
        74527 => X"62",  -- 98
        74528 => X"4E",  -- 78
        74529 => X"55",  -- 85
        74530 => X"58",  -- 88
        74531 => X"50",  -- 80
        74532 => X"3F",  -- 63
        74533 => X"2F",  -- 47
        74534 => X"29",  -- 41
        74535 => X"2B",  -- 43
        74536 => X"36",  -- 54
        74537 => X"3C",  -- 60
        74538 => X"3F",  -- 63
        74539 => X"42",  -- 66
        74540 => X"4C",  -- 76
        74541 => X"5A",  -- 90
        74542 => X"64",  -- 100
        74543 => X"63",  -- 99
        74544 => X"38",  -- 56
        74545 => X"3B",  -- 59
        74546 => X"47",  -- 71
        74547 => X"56",  -- 86
        74548 => X"62",  -- 98
        74549 => X"6C",  -- 108
        74550 => X"6B",  -- 107
        74551 => X"5E",  -- 94
        74552 => X"63",  -- 99
        74553 => X"71",  -- 113
        74554 => X"64",  -- 100
        74555 => X"57",  -- 87
        74556 => X"5A",  -- 90
        74557 => X"66",  -- 102
        74558 => X"7D",  -- 125
        74559 => X"87",  -- 135
        74560 => X"56",  -- 86
        74561 => X"55",  -- 85
        74562 => X"5B",  -- 91
        74563 => X"5D",  -- 93
        74564 => X"57",  -- 87
        74565 => X"59",  -- 89
        74566 => X"5F",  -- 95
        74567 => X"5D",  -- 93
        74568 => X"69",  -- 105
        74569 => X"60",  -- 96
        74570 => X"5B",  -- 91
        74571 => X"5C",  -- 92
        74572 => X"59",  -- 89
        74573 => X"53",  -- 83
        74574 => X"52",  -- 82
        74575 => X"56",  -- 86
        74576 => X"5A",  -- 90
        74577 => X"5D",  -- 93
        74578 => X"5A",  -- 90
        74579 => X"58",  -- 88
        74580 => X"5C",  -- 92
        74581 => X"56",  -- 86
        74582 => X"4C",  -- 76
        74583 => X"4B",  -- 75
        74584 => X"46",  -- 70
        74585 => X"4A",  -- 74
        74586 => X"5E",  -- 94
        74587 => X"5D",  -- 93
        74588 => X"50",  -- 80
        74589 => X"43",  -- 67
        74590 => X"49",  -- 73
        74591 => X"4E",  -- 78
        74592 => X"57",  -- 87
        74593 => X"41",  -- 65
        74594 => X"32",  -- 50
        74595 => X"34",  -- 52
        74596 => X"36",  -- 54
        74597 => X"34",  -- 52
        74598 => X"36",  -- 54
        74599 => X"3D",  -- 61
        74600 => X"2F",  -- 47
        74601 => X"29",  -- 41
        74602 => X"2C",  -- 44
        74603 => X"26",  -- 38
        74604 => X"4B",  -- 75
        74605 => X"2C",  -- 44
        74606 => X"23",  -- 35
        74607 => X"23",  -- 35
        74608 => X"2B",  -- 43
        74609 => X"50",  -- 80
        74610 => X"51",  -- 81
        74611 => X"3F",  -- 63
        74612 => X"3F",  -- 63
        74613 => X"3B",  -- 59
        74614 => X"3A",  -- 58
        74615 => X"31",  -- 49
        74616 => X"25",  -- 37
        74617 => X"26",  -- 38
        74618 => X"25",  -- 37
        74619 => X"27",  -- 39
        74620 => X"28",  -- 40
        74621 => X"20",  -- 32
        74622 => X"20",  -- 32
        74623 => X"2E",  -- 46
        74624 => X"3C",  -- 60
        74625 => X"3F",  -- 63
        74626 => X"3D",  -- 61
        74627 => X"3C",  -- 60
        74628 => X"3A",  -- 58
        74629 => X"2C",  -- 44
        74630 => X"20",  -- 32
        74631 => X"22",  -- 34
        74632 => X"34",  -- 52
        74633 => X"4B",  -- 75
        74634 => X"47",  -- 71
        74635 => X"3C",  -- 60
        74636 => X"42",  -- 66
        74637 => X"39",  -- 57
        74638 => X"25",  -- 37
        74639 => X"23",  -- 35
        74640 => X"21",  -- 33
        74641 => X"29",  -- 41
        74642 => X"33",  -- 51
        74643 => X"38",  -- 56
        74644 => X"35",  -- 53
        74645 => X"32",  -- 50
        74646 => X"34",  -- 52
        74647 => X"39",  -- 57
        74648 => X"2B",  -- 43
        74649 => X"29",  -- 41
        74650 => X"20",  -- 32
        74651 => X"1D",  -- 29
        74652 => X"24",  -- 36
        74653 => X"22",  -- 34
        74654 => X"1D",  -- 29
        74655 => X"1F",  -- 31
        74656 => X"17",  -- 23
        74657 => X"20",  -- 32
        74658 => X"28",  -- 40
        74659 => X"1F",  -- 31
        74660 => X"24",  -- 36
        74661 => X"2F",  -- 47
        74662 => X"2C",  -- 44
        74663 => X"36",  -- 54
        74664 => X"3F",  -- 63
        74665 => X"38",  -- 56
        74666 => X"28",  -- 40
        74667 => X"1D",  -- 29
        74668 => X"1C",  -- 28
        74669 => X"1B",  -- 27
        74670 => X"1A",  -- 26
        74671 => X"1D",  -- 29
        74672 => X"18",  -- 24
        74673 => X"1F",  -- 31
        74674 => X"23",  -- 35
        74675 => X"2A",  -- 42
        74676 => X"32",  -- 50
        74677 => X"30",  -- 48
        74678 => X"30",  -- 48
        74679 => X"3A",  -- 58
        74680 => X"34",  -- 52
        74681 => X"2F",  -- 47
        74682 => X"2D",  -- 45
        74683 => X"2F",  -- 47
        74684 => X"2B",  -- 43
        74685 => X"25",  -- 37
        74686 => X"28",  -- 40
        74687 => X"31",  -- 49
        74688 => X"36",  -- 54
        74689 => X"33",  -- 51
        74690 => X"2F",  -- 47
        74691 => X"2F",  -- 47
        74692 => X"2F",  -- 47
        74693 => X"2F",  -- 47
        74694 => X"2D",  -- 45
        74695 => X"2A",  -- 42
        74696 => X"26",  -- 38
        74697 => X"33",  -- 51
        74698 => X"3D",  -- 61
        74699 => X"3C",  -- 60
        74700 => X"40",  -- 64
        74701 => X"48",  -- 72
        74702 => X"4F",  -- 79
        74703 => X"4E",  -- 78
        74704 => X"53",  -- 83
        74705 => X"53",  -- 83
        74706 => X"5C",  -- 92
        74707 => X"5B",  -- 91
        74708 => X"55",  -- 85
        74709 => X"5E",  -- 94
        74710 => X"60",  -- 96
        74711 => X"4E",  -- 78
        74712 => X"4B",  -- 75
        74713 => X"49",  -- 73
        74714 => X"38",  -- 56
        74715 => X"32",  -- 50
        74716 => X"3C",  -- 60
        74717 => X"37",  -- 55
        74718 => X"28",  -- 40
        74719 => X"27",  -- 39
        74720 => X"40",  -- 64
        74721 => X"3C",  -- 60
        74722 => X"35",  -- 53
        74723 => X"34",  -- 52
        74724 => X"3B",  -- 59
        74725 => X"43",  -- 67
        74726 => X"3F",  -- 63
        74727 => X"37",  -- 55
        74728 => X"45",  -- 69
        74729 => X"3B",  -- 59
        74730 => X"37",  -- 55
        74731 => X"38",  -- 56
        74732 => X"3E",  -- 62
        74733 => X"4C",  -- 76
        74734 => X"4C",  -- 76
        74735 => X"3C",  -- 60
        74736 => X"35",  -- 53
        74737 => X"37",  -- 55
        74738 => X"37",  -- 55
        74739 => X"3F",  -- 63
        74740 => X"53",  -- 83
        74741 => X"63",  -- 99
        74742 => X"6B",  -- 107
        74743 => X"74",  -- 116
        74744 => X"6A",  -- 106
        74745 => X"5F",  -- 95
        74746 => X"53",  -- 83
        74747 => X"4C",  -- 76
        74748 => X"4E",  -- 78
        74749 => X"4D",  -- 77
        74750 => X"3D",  -- 61
        74751 => X"2D",  -- 45
        74752 => X"3A",  -- 58
        74753 => X"3A",  -- 58
        74754 => X"3E",  -- 62
        74755 => X"43",  -- 67
        74756 => X"49",  -- 73
        74757 => X"4E",  -- 78
        74758 => X"52",  -- 82
        74759 => X"54",  -- 84
        74760 => X"4D",  -- 77
        74761 => X"51",  -- 81
        74762 => X"54",  -- 84
        74763 => X"59",  -- 89
        74764 => X"5C",  -- 92
        74765 => X"60",  -- 96
        74766 => X"67",  -- 103
        74767 => X"6D",  -- 109
        74768 => X"64",  -- 100
        74769 => X"5A",  -- 90
        74770 => X"56",  -- 86
        74771 => X"56",  -- 86
        74772 => X"52",  -- 82
        74773 => X"49",  -- 73
        74774 => X"4C",  -- 76
        74775 => X"57",  -- 87
        74776 => X"4F",  -- 79
        74777 => X"41",  -- 65
        74778 => X"4C",  -- 76
        74779 => X"4B",  -- 75
        74780 => X"3D",  -- 61
        74781 => X"3F",  -- 63
        74782 => X"46",  -- 70
        74783 => X"4E",  -- 78
        74784 => X"3C",  -- 60
        74785 => X"42",  -- 66
        74786 => X"49",  -- 73
        74787 => X"4B",  -- 75
        74788 => X"47",  -- 71
        74789 => X"44",  -- 68
        74790 => X"44",  -- 68
        74791 => X"46",  -- 70
        74792 => X"44",  -- 68
        74793 => X"47",  -- 71
        74794 => X"4F",  -- 79
        74795 => X"54",  -- 84
        74796 => X"4F",  -- 79
        74797 => X"48",  -- 72
        74798 => X"49",  -- 73
        74799 => X"4F",  -- 79
        74800 => X"61",  -- 97
        74801 => X"5D",  -- 93
        74802 => X"4E",  -- 78
        74803 => X"45",  -- 69
        74804 => X"47",  -- 71
        74805 => X"45",  -- 69
        74806 => X"42",  -- 66
        74807 => X"47",  -- 71
        74808 => X"48",  -- 72
        74809 => X"3D",  -- 61
        74810 => X"51",  -- 81
        74811 => X"55",  -- 85
        74812 => X"6A",  -- 106
        74813 => X"62",  -- 98
        74814 => X"59",  -- 89
        74815 => X"57",  -- 87
        74816 => X"6A",  -- 106
        74817 => X"75",  -- 117
        74818 => X"61",  -- 97
        74819 => X"61",  -- 97
        74820 => X"64",  -- 100
        74821 => X"5D",  -- 93
        74822 => X"64",  -- 100
        74823 => X"58",  -- 88
        74824 => X"4B",  -- 75
        74825 => X"44",  -- 68
        74826 => X"66",  -- 102
        74827 => X"6B",  -- 107
        74828 => X"5E",  -- 94
        74829 => X"4D",  -- 77
        74830 => X"66",  -- 102
        74831 => X"6A",  -- 106
        74832 => X"41",  -- 65
        74833 => X"49",  -- 73
        74834 => X"70",  -- 112
        74835 => X"7D",  -- 125
        74836 => X"9A",  -- 154
        74837 => X"91",  -- 145
        74838 => X"93",  -- 147
        74839 => X"8D",  -- 141
        74840 => X"92",  -- 146
        74841 => X"90",  -- 144
        74842 => X"83",  -- 131
        74843 => X"7E",  -- 126
        74844 => X"6D",  -- 109
        74845 => X"3B",  -- 59
        74846 => X"41",  -- 65
        74847 => X"38",  -- 56
        74848 => X"4F",  -- 79
        74849 => X"41",  -- 65
        74850 => X"3B",  -- 59
        74851 => X"41",  -- 65
        74852 => X"44",  -- 68
        74853 => X"3F",  -- 63
        74854 => X"3C",  -- 60
        74855 => X"3F",  -- 63
        74856 => X"37",  -- 55
        74857 => X"34",  -- 52
        74858 => X"35",  -- 53
        74859 => X"38",  -- 56
        74860 => X"31",  -- 49
        74861 => X"22",  -- 34
        74862 => X"19",  -- 25
        74863 => X"17",  -- 23
        74864 => X"1B",  -- 27
        74865 => X"27",  -- 39
        74866 => X"36",  -- 54
        74867 => X"38",  -- 56
        74868 => X"32",  -- 50
        74869 => X"3A",  -- 58
        74870 => X"4D",  -- 77
        74871 => X"55",  -- 85
        74872 => X"50",  -- 80
        74873 => X"4B",  -- 75
        74874 => X"4E",  -- 78
        74875 => X"59",  -- 89
        74876 => X"5F",  -- 95
        74877 => X"57",  -- 87
        74878 => X"5B",  -- 91
        74879 => X"74",  -- 116
        74880 => X"67",  -- 103
        74881 => X"61",  -- 97
        74882 => X"61",  -- 97
        74883 => X"61",  -- 97
        74884 => X"5D",  -- 93
        74885 => X"60",  -- 96
        74886 => X"63",  -- 99
        74887 => X"5F",  -- 95
        74888 => X"63",  -- 99
        74889 => X"61",  -- 97
        74890 => X"5D",  -- 93
        74891 => X"57",  -- 87
        74892 => X"55",  -- 85
        74893 => X"57",  -- 87
        74894 => X"5B",  -- 91
        74895 => X"5F",  -- 95
        74896 => X"65",  -- 101
        74897 => X"64",  -- 100
        74898 => X"5B",  -- 91
        74899 => X"58",  -- 88
        74900 => X"5E",  -- 94
        74901 => X"5C",  -- 92
        74902 => X"55",  -- 85
        74903 => X"57",  -- 87
        74904 => X"5F",  -- 95
        74905 => X"51",  -- 81
        74906 => X"65",  -- 101
        74907 => X"46",  -- 70
        74908 => X"46",  -- 70
        74909 => X"49",  -- 73
        74910 => X"55",  -- 85
        74911 => X"5B",  -- 91
        74912 => X"5D",  -- 93
        74913 => X"41",  -- 65
        74914 => X"2D",  -- 45
        74915 => X"34",  -- 52
        74916 => X"41",  -- 65
        74917 => X"40",  -- 64
        74918 => X"31",  -- 49
        74919 => X"27",  -- 39
        74920 => X"29",  -- 41
        74921 => X"25",  -- 37
        74922 => X"2B",  -- 43
        74923 => X"2A",  -- 42
        74924 => X"4C",  -- 76
        74925 => X"35",  -- 53
        74926 => X"2E",  -- 46
        74927 => X"2F",  -- 47
        74928 => X"3A",  -- 58
        74929 => X"4D",  -- 77
        74930 => X"62",  -- 98
        74931 => X"40",  -- 64
        74932 => X"42",  -- 66
        74933 => X"41",  -- 65
        74934 => X"40",  -- 64
        74935 => X"2E",  -- 46
        74936 => X"2A",  -- 42
        74937 => X"24",  -- 36
        74938 => X"1E",  -- 30
        74939 => X"24",  -- 36
        74940 => X"2B",  -- 43
        74941 => X"24",  -- 36
        74942 => X"22",  -- 34
        74943 => X"2E",  -- 46
        74944 => X"42",  -- 66
        74945 => X"43",  -- 67
        74946 => X"43",  -- 67
        74947 => X"46",  -- 70
        74948 => X"42",  -- 66
        74949 => X"2F",  -- 47
        74950 => X"24",  -- 36
        74951 => X"2C",  -- 44
        74952 => X"3A",  -- 58
        74953 => X"44",  -- 68
        74954 => X"3D",  -- 61
        74955 => X"38",  -- 56
        74956 => X"42",  -- 66
        74957 => X"39",  -- 57
        74958 => X"25",  -- 37
        74959 => X"21",  -- 33
        74960 => X"23",  -- 35
        74961 => X"2A",  -- 42
        74962 => X"35",  -- 53
        74963 => X"3C",  -- 60
        74964 => X"3C",  -- 60
        74965 => X"38",  -- 56
        74966 => X"39",  -- 57
        74967 => X"3E",  -- 62
        74968 => X"34",  -- 52
        74969 => X"2B",  -- 43
        74970 => X"1E",  -- 30
        74971 => X"1F",  -- 31
        74972 => X"27",  -- 39
        74973 => X"22",  -- 34
        74974 => X"1A",  -- 26
        74975 => X"1C",  -- 28
        74976 => X"15",  -- 21
        74977 => X"1D",  -- 29
        74978 => X"20",  -- 32
        74979 => X"18",  -- 24
        74980 => X"2E",  -- 46
        74981 => X"46",  -- 70
        74982 => X"34",  -- 52
        74983 => X"25",  -- 37
        74984 => X"3F",  -- 63
        74985 => X"2D",  -- 45
        74986 => X"1E",  -- 30
        74987 => X"1E",  -- 30
        74988 => X"22",  -- 34
        74989 => X"21",  -- 33
        74990 => X"1D",  -- 29
        74991 => X"1C",  -- 28
        74992 => X"1C",  -- 28
        74993 => X"21",  -- 33
        74994 => X"20",  -- 32
        74995 => X"23",  -- 35
        74996 => X"2A",  -- 42
        74997 => X"2D",  -- 45
        74998 => X"31",  -- 49
        74999 => X"3E",  -- 62
        75000 => X"2E",  -- 46
        75001 => X"2B",  -- 43
        75002 => X"2C",  -- 44
        75003 => X"2E",  -- 46
        75004 => X"2C",  -- 44
        75005 => X"27",  -- 39
        75006 => X"29",  -- 41
        75007 => X"2F",  -- 47
        75008 => X"31",  -- 49
        75009 => X"2F",  -- 47
        75010 => X"2C",  -- 44
        75011 => X"2D",  -- 45
        75012 => X"31",  -- 49
        75013 => X"33",  -- 51
        75014 => X"31",  -- 49
        75015 => X"30",  -- 48
        75016 => X"34",  -- 52
        75017 => X"3B",  -- 59
        75018 => X"43",  -- 67
        75019 => X"45",  -- 69
        75020 => X"47",  -- 71
        75021 => X"4D",  -- 77
        75022 => X"4C",  -- 76
        75023 => X"49",  -- 73
        75024 => X"4F",  -- 79
        75025 => X"4E",  -- 78
        75026 => X"4F",  -- 79
        75027 => X"49",  -- 73
        75028 => X"44",  -- 68
        75029 => X"4C",  -- 76
        75030 => X"4D",  -- 77
        75031 => X"3C",  -- 60
        75032 => X"3E",  -- 62
        75033 => X"38",  -- 56
        75034 => X"30",  -- 48
        75035 => X"37",  -- 55
        75036 => X"44",  -- 68
        75037 => X"41",  -- 65
        75038 => X"3A",  -- 58
        75039 => X"3D",  -- 61
        75040 => X"44",  -- 68
        75041 => X"3C",  -- 60
        75042 => X"35",  -- 53
        75043 => X"38",  -- 56
        75044 => X"3D",  -- 61
        75045 => X"3B",  -- 59
        75046 => X"38",  -- 56
        75047 => X"35",  -- 53
        75048 => X"39",  -- 57
        75049 => X"37",  -- 55
        75050 => X"38",  -- 56
        75051 => X"34",  -- 52
        75052 => X"31",  -- 49
        75053 => X"3D",  -- 61
        75054 => X"48",  -- 72
        75055 => X"47",  -- 71
        75056 => X"3C",  -- 60
        75057 => X"47",  -- 71
        75058 => X"4A",  -- 74
        75059 => X"4B",  -- 75
        75060 => X"4F",  -- 79
        75061 => X"55",  -- 85
        75062 => X"5E",  -- 94
        75063 => X"6D",  -- 109
        75064 => X"67",  -- 103
        75065 => X"6E",  -- 110
        75066 => X"66",  -- 102
        75067 => X"4F",  -- 79
        75068 => X"44",  -- 68
        75069 => X"47",  -- 71
        75070 => X"48",  -- 72
        75071 => X"41",  -- 65
        75072 => X"3E",  -- 62
        75073 => X"3E",  -- 62
        75074 => X"3B",  -- 59
        75075 => X"3D",  -- 61
        75076 => X"43",  -- 67
        75077 => X"4C",  -- 76
        75078 => X"53",  -- 83
        75079 => X"57",  -- 87
        75080 => X"5C",  -- 92
        75081 => X"59",  -- 89
        75082 => X"56",  -- 86
        75083 => X"56",  -- 86
        75084 => X"5A",  -- 90
        75085 => X"63",  -- 99
        75086 => X"6C",  -- 108
        75087 => X"71",  -- 113
        75088 => X"63",  -- 99
        75089 => X"5A",  -- 90
        75090 => X"54",  -- 84
        75091 => X"55",  -- 85
        75092 => X"58",  -- 88
        75093 => X"53",  -- 83
        75094 => X"4C",  -- 76
        75095 => X"45",  -- 69
        75096 => X"46",  -- 70
        75097 => X"44",  -- 68
        75098 => X"43",  -- 67
        75099 => X"4B",  -- 75
        75100 => X"47",  -- 71
        75101 => X"47",  -- 71
        75102 => X"50",  -- 80
        75103 => X"49",  -- 73
        75104 => X"40",  -- 64
        75105 => X"44",  -- 68
        75106 => X"48",  -- 72
        75107 => X"49",  -- 73
        75108 => X"45",  -- 69
        75109 => X"42",  -- 66
        75110 => X"43",  -- 67
        75111 => X"46",  -- 70
        75112 => X"44",  -- 68
        75113 => X"44",  -- 68
        75114 => X"4A",  -- 74
        75115 => X"51",  -- 81
        75116 => X"4C",  -- 76
        75117 => X"43",  -- 67
        75118 => X"43",  -- 67
        75119 => X"4A",  -- 74
        75120 => X"41",  -- 65
        75121 => X"49",  -- 73
        75122 => X"49",  -- 73
        75123 => X"48",  -- 72
        75124 => X"4C",  -- 76
        75125 => X"4A",  -- 74
        75126 => X"45",  -- 69
        75127 => X"48",  -- 72
        75128 => X"47",  -- 71
        75129 => X"53",  -- 83
        75130 => X"61",  -- 97
        75131 => X"4C",  -- 76
        75132 => X"59",  -- 89
        75133 => X"6A",  -- 106
        75134 => X"60",  -- 96
        75135 => X"48",  -- 72
        75136 => X"50",  -- 80
        75137 => X"7C",  -- 124
        75138 => X"62",  -- 98
        75139 => X"5F",  -- 95
        75140 => X"67",  -- 103
        75141 => X"57",  -- 87
        75142 => X"61",  -- 97
        75143 => X"5A",  -- 90
        75144 => X"5E",  -- 94
        75145 => X"55",  -- 85
        75146 => X"69",  -- 105
        75147 => X"5F",  -- 95
        75148 => X"5D",  -- 93
        75149 => X"51",  -- 81
        75150 => X"5C",  -- 92
        75151 => X"48",  -- 72
        75152 => X"2D",  -- 45
        75153 => X"40",  -- 64
        75154 => X"62",  -- 98
        75155 => X"7F",  -- 127
        75156 => X"9A",  -- 154
        75157 => X"9A",  -- 154
        75158 => X"94",  -- 148
        75159 => X"87",  -- 135
        75160 => X"99",  -- 153
        75161 => X"87",  -- 135
        75162 => X"85",  -- 133
        75163 => X"85",  -- 133
        75164 => X"74",  -- 116
        75165 => X"42",  -- 66
        75166 => X"33",  -- 51
        75167 => X"39",  -- 57
        75168 => X"3F",  -- 63
        75169 => X"43",  -- 67
        75170 => X"51",  -- 81
        75171 => X"5D",  -- 93
        75172 => X"4D",  -- 77
        75173 => X"35",  -- 53
        75174 => X"32",  -- 50
        75175 => X"42",  -- 66
        75176 => X"26",  -- 38
        75177 => X"2A",  -- 42
        75178 => X"2F",  -- 47
        75179 => X"2B",  -- 43
        75180 => X"1B",  -- 27
        75181 => X"10",  -- 16
        75182 => X"14",  -- 20
        75183 => X"22",  -- 34
        75184 => X"48",  -- 72
        75185 => X"42",  -- 66
        75186 => X"3D",  -- 61
        75187 => X"3A",  -- 58
        75188 => X"3C",  -- 60
        75189 => X"4F",  -- 79
        75190 => X"64",  -- 100
        75191 => X"69",  -- 105
        75192 => X"6D",  -- 109
        75193 => X"5A",  -- 90
        75194 => X"56",  -- 86
        75195 => X"53",  -- 83
        75196 => X"66",  -- 102
        75197 => X"6D",  -- 109
        75198 => X"4D",  -- 77
        75199 => X"48",  -- 72
        75200 => X"66",  -- 102
        75201 => X"5F",  -- 95
        75202 => X"60",  -- 96
        75203 => X"63",  -- 99
        75204 => X"61",  -- 97
        75205 => X"61",  -- 97
        75206 => X"5D",  -- 93
        75207 => X"53",  -- 83
        75208 => X"4A",  -- 74
        75209 => X"4F",  -- 79
        75210 => X"51",  -- 81
        75211 => X"4C",  -- 76
        75212 => X"4D",  -- 77
        75213 => X"58",  -- 88
        75214 => X"61",  -- 97
        75215 => X"63",  -- 99
        75216 => X"63",  -- 99
        75217 => X"60",  -- 96
        75218 => X"55",  -- 85
        75219 => X"51",  -- 81
        75220 => X"5A",  -- 90
        75221 => X"5D",  -- 93
        75222 => X"5C",  -- 92
        75223 => X"60",  -- 96
        75224 => X"66",  -- 102
        75225 => X"4E",  -- 78
        75226 => X"62",  -- 98
        75227 => X"2F",  -- 47
        75228 => X"37",  -- 55
        75229 => X"47",  -- 71
        75230 => X"58",  -- 88
        75231 => X"60",  -- 96
        75232 => X"54",  -- 84
        75233 => X"47",  -- 71
        75234 => X"3D",  -- 61
        75235 => X"3E",  -- 62
        75236 => X"3E",  -- 62
        75237 => X"35",  -- 53
        75238 => X"2A",  -- 42
        75239 => X"24",  -- 36
        75240 => X"33",  -- 51
        75241 => X"2C",  -- 44
        75242 => X"2F",  -- 47
        75243 => X"30",  -- 48
        75244 => X"4C",  -- 76
        75245 => X"40",  -- 64
        75246 => X"40",  -- 64
        75247 => X"42",  -- 66
        75248 => X"41",  -- 65
        75249 => X"40",  -- 64
        75250 => X"58",  -- 88
        75251 => X"40",  -- 64
        75252 => X"3E",  -- 62
        75253 => X"42",  -- 66
        75254 => X"31",  -- 49
        75255 => X"20",  -- 32
        75256 => X"29",  -- 41
        75257 => X"27",  -- 39
        75258 => X"1E",  -- 30
        75259 => X"1C",  -- 28
        75260 => X"25",  -- 37
        75261 => X"27",  -- 39
        75262 => X"28",  -- 40
        75263 => X"2E",  -- 46
        75264 => X"43",  -- 67
        75265 => X"40",  -- 64
        75266 => X"40",  -- 64
        75267 => X"47",  -- 71
        75268 => X"44",  -- 68
        75269 => X"2E",  -- 46
        75270 => X"20",  -- 32
        75271 => X"29",  -- 41
        75272 => X"3A",  -- 58
        75273 => X"3E",  -- 62
        75274 => X"38",  -- 56
        75275 => X"38",  -- 56
        75276 => X"3E",  -- 62
        75277 => X"33",  -- 51
        75278 => X"21",  -- 33
        75279 => X"1B",  -- 27
        75280 => X"1B",  -- 27
        75281 => X"28",  -- 40
        75282 => X"33",  -- 51
        75283 => X"35",  -- 53
        75284 => X"34",  -- 52
        75285 => X"34",  -- 52
        75286 => X"32",  -- 50
        75287 => X"2F",  -- 47
        75288 => X"2E",  -- 46
        75289 => X"28",  -- 40
        75290 => X"20",  -- 32
        75291 => X"26",  -- 38
        75292 => X"2E",  -- 46
        75293 => X"25",  -- 37
        75294 => X"19",  -- 25
        75295 => X"1A",  -- 26
        75296 => X"16",  -- 22
        75297 => X"1D",  -- 29
        75298 => X"1F",  -- 31
        75299 => X"16",  -- 22
        75300 => X"2C",  -- 44
        75301 => X"44",  -- 68
        75302 => X"36",  -- 54
        75303 => X"2B",  -- 43
        75304 => X"3C",  -- 60
        75305 => X"28",  -- 40
        75306 => X"23",  -- 35
        75307 => X"2D",  -- 45
        75308 => X"2F",  -- 47
        75309 => X"28",  -- 40
        75310 => X"1F",  -- 31
        75311 => X"19",  -- 25
        75312 => X"28",  -- 40
        75313 => X"29",  -- 41
        75314 => X"21",  -- 33
        75315 => X"1F",  -- 31
        75316 => X"28",  -- 40
        75317 => X"2C",  -- 44
        75318 => X"2F",  -- 47
        75319 => X"37",  -- 55
        75320 => X"2B",  -- 43
        75321 => X"2A",  -- 42
        75322 => X"2D",  -- 45
        75323 => X"30",  -- 48
        75324 => X"30",  -- 48
        75325 => X"2D",  -- 45
        75326 => X"2F",  -- 47
        75327 => X"34",  -- 52
        75328 => X"34",  -- 52
        75329 => X"31",  -- 49
        75330 => X"30",  -- 48
        75331 => X"31",  -- 49
        75332 => X"35",  -- 53
        75333 => X"3A",  -- 58
        75334 => X"3C",  -- 60
        75335 => X"3C",  -- 60
        75336 => X"3D",  -- 61
        75337 => X"41",  -- 65
        75338 => X"45",  -- 69
        75339 => X"47",  -- 71
        75340 => X"49",  -- 73
        75341 => X"49",  -- 73
        75342 => X"49",  -- 73
        75343 => X"46",  -- 70
        75344 => X"46",  -- 70
        75345 => X"3F",  -- 63
        75346 => X"3B",  -- 59
        75347 => X"38",  -- 56
        75348 => X"35",  -- 53
        75349 => X"34",  -- 52
        75350 => X"35",  -- 53
        75351 => X"32",  -- 50
        75352 => X"33",  -- 51
        75353 => X"35",  -- 53
        75354 => X"3B",  -- 59
        75355 => X"45",  -- 69
        75356 => X"47",  -- 71
        75357 => X"3D",  -- 61
        75358 => X"3C",  -- 60
        75359 => X"47",  -- 71
        75360 => X"44",  -- 68
        75361 => X"37",  -- 55
        75362 => X"35",  -- 53
        75363 => X"3E",  -- 62
        75364 => X"42",  -- 66
        75365 => X"3B",  -- 59
        75366 => X"36",  -- 54
        75367 => X"3B",  -- 59
        75368 => X"30",  -- 48
        75369 => X"34",  -- 52
        75370 => X"3B",  -- 59
        75371 => X"37",  -- 55
        75372 => X"30",  -- 48
        75373 => X"39",  -- 57
        75374 => X"49",  -- 73
        75375 => X"4D",  -- 77
        75376 => X"44",  -- 68
        75377 => X"53",  -- 83
        75378 => X"5A",  -- 90
        75379 => X"56",  -- 86
        75380 => X"50",  -- 80
        75381 => X"4B",  -- 75
        75382 => X"50",  -- 80
        75383 => X"5F",  -- 95
        75384 => X"63",  -- 99
        75385 => X"60",  -- 96
        75386 => X"5D",  -- 93
        75387 => X"57",  -- 87
        75388 => X"4C",  -- 76
        75389 => X"42",  -- 66
        75390 => X"4C",  -- 76
        75391 => X"5E",  -- 94
        75392 => X"3D",  -- 61
        75393 => X"40",  -- 64
        75394 => X"41",  -- 65
        75395 => X"3E",  -- 62
        75396 => X"42",  -- 66
        75397 => X"4C",  -- 76
        75398 => X"58",  -- 88
        75399 => X"5E",  -- 94
        75400 => X"61",  -- 97
        75401 => X"59",  -- 89
        75402 => X"52",  -- 82
        75403 => X"4F",  -- 79
        75404 => X"53",  -- 83
        75405 => X"5C",  -- 92
        75406 => X"66",  -- 102
        75407 => X"6C",  -- 108
        75408 => X"69",  -- 105
        75409 => X"5E",  -- 94
        75410 => X"54",  -- 84
        75411 => X"54",  -- 84
        75412 => X"5C",  -- 92
        75413 => X"59",  -- 89
        75414 => X"46",  -- 70
        75415 => X"33",  -- 51
        75416 => X"3D",  -- 61
        75417 => X"44",  -- 68
        75418 => X"3C",  -- 60
        75419 => X"49",  -- 73
        75420 => X"4C",  -- 76
        75421 => X"46",  -- 70
        75422 => X"51",  -- 81
        75423 => X"42",  -- 66
        75424 => X"4A",  -- 74
        75425 => X"4B",  -- 75
        75426 => X"4C",  -- 76
        75427 => X"49",  -- 73
        75428 => X"45",  -- 69
        75429 => X"42",  -- 66
        75430 => X"42",  -- 66
        75431 => X"44",  -- 68
        75432 => X"49",  -- 73
        75433 => X"43",  -- 67
        75434 => X"42",  -- 66
        75435 => X"46",  -- 70
        75436 => X"4B",  -- 75
        75437 => X"4C",  -- 76
        75438 => X"49",  -- 73
        75439 => X"44",  -- 68
        75440 => X"44",  -- 68
        75441 => X"4D",  -- 77
        75442 => X"4E",  -- 78
        75443 => X"4C",  -- 76
        75444 => X"4D",  -- 77
        75445 => X"47",  -- 71
        75446 => X"3C",  -- 60
        75447 => X"39",  -- 57
        75448 => X"45",  -- 69
        75449 => X"4D",  -- 77
        75450 => X"58",  -- 88
        75451 => X"48",  -- 72
        75452 => X"4A",  -- 74
        75453 => X"57",  -- 87
        75454 => X"51",  -- 81
        75455 => X"48",  -- 72
        75456 => X"63",  -- 99
        75457 => X"7D",  -- 125
        75458 => X"71",  -- 113
        75459 => X"6A",  -- 106
        75460 => X"69",  -- 105
        75461 => X"5D",  -- 93
        75462 => X"5E",  -- 94
        75463 => X"5A",  -- 90
        75464 => X"5C",  -- 92
        75465 => X"56",  -- 86
        75466 => X"53",  -- 83
        75467 => X"53",  -- 83
        75468 => X"45",  -- 69
        75469 => X"4B",  -- 75
        75470 => X"46",  -- 70
        75471 => X"3A",  -- 58
        75472 => X"3A",  -- 58
        75473 => X"4C",  -- 76
        75474 => X"66",  -- 102
        75475 => X"8F",  -- 143
        75476 => X"97",  -- 151
        75477 => X"8B",  -- 139
        75478 => X"85",  -- 133
        75479 => X"85",  -- 133
        75480 => X"8A",  -- 138
        75481 => X"74",  -- 116
        75482 => X"7D",  -- 125
        75483 => X"7A",  -- 122
        75484 => X"6C",  -- 108
        75485 => X"4E",  -- 78
        75486 => X"34",  -- 52
        75487 => X"40",  -- 64
        75488 => X"30",  -- 48
        75489 => X"2E",  -- 46
        75490 => X"36",  -- 54
        75491 => X"42",  -- 66
        75492 => X"3E",  -- 62
        75493 => X"29",  -- 41
        75494 => X"14",  -- 20
        75495 => X"0C",  -- 12
        75496 => X"0F",  -- 15
        75497 => X"12",  -- 18
        75498 => X"17",  -- 23
        75499 => X"1A",  -- 26
        75500 => X"22",  -- 34
        75501 => X"2F",  -- 47
        75502 => X"41",  -- 65
        75503 => X"4F",  -- 79
        75504 => X"50",  -- 80
        75505 => X"50",  -- 80
        75506 => X"5C",  -- 92
        75507 => X"6D",  -- 109
        75508 => X"79",  -- 121
        75509 => X"7D",  -- 125
        75510 => X"6F",  -- 111
        75511 => X"58",  -- 88
        75512 => X"4A",  -- 74
        75513 => X"3A",  -- 58
        75514 => X"43",  -- 67
        75515 => X"3C",  -- 60
        75516 => X"53",  -- 83
        75517 => X"63",  -- 99
        75518 => X"36",  -- 54
        75519 => X"2A",  -- 42
        75520 => X"60",  -- 96
        75521 => X"58",  -- 88
        75522 => X"59",  -- 89
        75523 => X"5E",  -- 94
        75524 => X"60",  -- 96
        75525 => X"62",  -- 98
        75526 => X"5F",  -- 95
        75527 => X"54",  -- 84
        75528 => X"37",  -- 55
        75529 => X"3D",  -- 61
        75530 => X"3E",  -- 62
        75531 => X"38",  -- 56
        75532 => X"3C",  -- 60
        75533 => X"4C",  -- 76
        75534 => X"59",  -- 89
        75535 => X"5C",  -- 92
        75536 => X"58",  -- 88
        75537 => X"59",  -- 89
        75538 => X"54",  -- 84
        75539 => X"54",  -- 84
        75540 => X"5F",  -- 95
        75541 => X"62",  -- 98
        75542 => X"5F",  -- 95
        75543 => X"62",  -- 98
        75544 => X"62",  -- 98
        75545 => X"4D",  -- 77
        75546 => X"61",  -- 97
        75547 => X"2B",  -- 43
        75548 => X"32",  -- 50
        75549 => X"46",  -- 70
        75550 => X"59",  -- 89
        75551 => X"60",  -- 96
        75552 => X"56",  -- 86
        75553 => X"58",  -- 88
        75554 => X"56",  -- 86
        75555 => X"4A",  -- 74
        75556 => X"37",  -- 55
        75557 => X"26",  -- 38
        75558 => X"22",  -- 34
        75559 => X"24",  -- 36
        75560 => X"39",  -- 57
        75561 => X"33",  -- 51
        75562 => X"36",  -- 54
        75563 => X"3A",  -- 58
        75564 => X"4E",  -- 78
        75565 => X"48",  -- 72
        75566 => X"49",  -- 73
        75567 => X"49",  -- 73
        75568 => X"44",  -- 68
        75569 => X"40",  -- 64
        75570 => X"51",  -- 81
        75571 => X"52",  -- 82
        75572 => X"3E",  -- 62
        75573 => X"40",  -- 64
        75574 => X"24",  -- 36
        75575 => X"24",  -- 36
        75576 => X"25",  -- 37
        75577 => X"2F",  -- 47
        75578 => X"23",  -- 35
        75579 => X"11",  -- 17
        75580 => X"16",  -- 22
        75581 => X"25",  -- 37
        75582 => X"2A",  -- 42
        75583 => X"2A",  -- 42
        75584 => X"48",  -- 72
        75585 => X"44",  -- 68
        75586 => X"42",  -- 66
        75587 => X"49",  -- 73
        75588 => X"48",  -- 72
        75589 => X"31",  -- 49
        75590 => X"20",  -- 32
        75591 => X"25",  -- 37
        75592 => X"35",  -- 53
        75593 => X"39",  -- 57
        75594 => X"3B",  -- 59
        75595 => X"3D",  -- 61
        75596 => X"3E",  -- 62
        75597 => X"33",  -- 51
        75598 => X"24",  -- 36
        75599 => X"1D",  -- 29
        75600 => X"1C",  -- 28
        75601 => X"30",  -- 48
        75602 => X"3B",  -- 59
        75603 => X"34",  -- 52
        75604 => X"32",  -- 50
        75605 => X"39",  -- 57
        75606 => X"34",  -- 52
        75607 => X"26",  -- 38
        75608 => X"22",  -- 34
        75609 => X"24",  -- 36
        75610 => X"26",  -- 38
        75611 => X"2F",  -- 47
        75612 => X"36",  -- 54
        75613 => X"2A",  -- 42
        75614 => X"1C",  -- 28
        75615 => X"1C",  -- 28
        75616 => X"13",  -- 19
        75617 => X"1B",  -- 27
        75618 => X"25",  -- 37
        75619 => X"21",  -- 33
        75620 => X"2A",  -- 42
        75621 => X"36",  -- 54
        75622 => X"33",  -- 51
        75623 => X"3F",  -- 63
        75624 => X"3A",  -- 58
        75625 => X"28",  -- 40
        75626 => X"2B",  -- 43
        75627 => X"37",  -- 55
        75628 => X"31",  -- 49
        75629 => X"27",  -- 39
        75630 => X"22",  -- 34
        75631 => X"1B",  -- 27
        75632 => X"33",  -- 51
        75633 => X"2F",  -- 47
        75634 => X"23",  -- 35
        75635 => X"1F",  -- 31
        75636 => X"2A",  -- 42
        75637 => X"30",  -- 48
        75638 => X"2D",  -- 45
        75639 => X"2F",  -- 47
        75640 => X"2E",  -- 46
        75641 => X"2F",  -- 47
        75642 => X"33",  -- 51
        75643 => X"36",  -- 54
        75644 => X"35",  -- 53
        75645 => X"33",  -- 51
        75646 => X"34",  -- 52
        75647 => X"37",  -- 55
        75648 => X"41",  -- 65
        75649 => X"3D",  -- 61
        75650 => X"37",  -- 55
        75651 => X"36",  -- 54
        75652 => X"39",  -- 57
        75653 => X"3D",  -- 61
        75654 => X"40",  -- 64
        75655 => X"41",  -- 65
        75656 => X"42",  -- 66
        75657 => X"43",  -- 67
        75658 => X"46",  -- 70
        75659 => X"48",  -- 72
        75660 => X"46",  -- 70
        75661 => X"44",  -- 68
        75662 => X"47",  -- 71
        75663 => X"4B",  -- 75
        75664 => X"39",  -- 57
        75665 => X"34",  -- 52
        75666 => X"35",  -- 53
        75667 => X"3A",  -- 58
        75668 => X"36",  -- 54
        75669 => X"26",  -- 38
        75670 => X"24",  -- 36
        75671 => X"31",  -- 49
        75672 => X"41",  -- 65
        75673 => X"3A",  -- 58
        75674 => X"3E",  -- 62
        75675 => X"43",  -- 67
        75676 => X"3B",  -- 59
        75677 => X"31",  -- 49
        75678 => X"36",  -- 54
        75679 => X"40",  -- 64
        75680 => X"41",  -- 65
        75681 => X"35",  -- 53
        75682 => X"38",  -- 56
        75683 => X"46",  -- 70
        75684 => X"4A",  -- 74
        75685 => X"3E",  -- 62
        75686 => X"3A",  -- 58
        75687 => X"42",  -- 66
        75688 => X"37",  -- 55
        75689 => X"31",  -- 49
        75690 => X"34",  -- 52
        75691 => X"39",  -- 57
        75692 => X"3D",  -- 61
        75693 => X"47",  -- 71
        75694 => X"49",  -- 73
        75695 => X"41",  -- 65
        75696 => X"44",  -- 68
        75697 => X"53",  -- 83
        75698 => X"59",  -- 89
        75699 => X"55",  -- 85
        75700 => X"50",  -- 80
        75701 => X"48",  -- 72
        75702 => X"46",  -- 70
        75703 => X"50",  -- 80
        75704 => X"67",  -- 103
        75705 => X"54",  -- 84
        75706 => X"4F",  -- 79
        75707 => X"5B",  -- 91
        75708 => X"5D",  -- 93
        75709 => X"4E",  -- 78
        75710 => X"47",  -- 71
        75711 => X"4B",  -- 75
        75712 => X"33",  -- 51
        75713 => X"3D",  -- 61
        75714 => X"43",  -- 67
        75715 => X"42",  -- 66
        75716 => X"45",  -- 69
        75717 => X"51",  -- 81
        75718 => X"61",  -- 97
        75719 => X"6A",  -- 106
        75720 => X"68",  -- 104
        75721 => X"61",  -- 97
        75722 => X"58",  -- 88
        75723 => X"54",  -- 84
        75724 => X"57",  -- 87
        75725 => X"5E",  -- 94
        75726 => X"67",  -- 103
        75727 => X"6C",  -- 108
        75728 => X"6C",  -- 108
        75729 => X"5E",  -- 94
        75730 => X"51",  -- 81
        75731 => X"4C",  -- 76
        75732 => X"52",  -- 82
        75733 => X"50",  -- 80
        75734 => X"39",  -- 57
        75735 => X"20",  -- 32
        75736 => X"2D",  -- 45
        75737 => X"42",  -- 66
        75738 => X"40",  -- 64
        75739 => X"49",  -- 73
        75740 => X"43",  -- 67
        75741 => X"34",  -- 52
        75742 => X"45",  -- 69
        75743 => X"46",  -- 70
        75744 => X"51",  -- 81
        75745 => X"50",  -- 80
        75746 => X"4E",  -- 78
        75747 => X"4B",  -- 75
        75748 => X"46",  -- 70
        75749 => X"44",  -- 68
        75750 => X"46",  -- 70
        75751 => X"47",  -- 71
        75752 => X"49",  -- 73
        75753 => X"48",  -- 72
        75754 => X"44",  -- 68
        75755 => X"40",  -- 64
        75756 => X"47",  -- 71
        75757 => X"50",  -- 80
        75758 => X"4D",  -- 77
        75759 => X"43",  -- 67
        75760 => X"50",  -- 80
        75761 => X"53",  -- 83
        75762 => X"49",  -- 73
        75763 => X"42",  -- 66
        75764 => X"48",  -- 72
        75765 => X"4B",  -- 75
        75766 => X"47",  -- 71
        75767 => X"47",  -- 71
        75768 => X"4A",  -- 74
        75769 => X"3D",  -- 61
        75770 => X"47",  -- 71
        75771 => X"50",  -- 80
        75772 => X"48",  -- 72
        75773 => X"3E",  -- 62
        75774 => X"3D",  -- 61
        75775 => X"59",  -- 89
        75776 => X"6A",  -- 106
        75777 => X"58",  -- 88
        75778 => X"66",  -- 102
        75779 => X"61",  -- 97
        75780 => X"56",  -- 86
        75781 => X"5B",  -- 91
        75782 => X"51",  -- 81
        75783 => X"4F",  -- 79
        75784 => X"5A",  -- 90
        75785 => X"52",  -- 82
        75786 => X"50",  -- 80
        75787 => X"4E",  -- 78
        75788 => X"44",  -- 68
        75789 => X"3C",  -- 60
        75790 => X"39",  -- 57
        75791 => X"36",  -- 54
        75792 => X"3B",  -- 59
        75793 => X"5B",  -- 91
        75794 => X"77",  -- 119
        75795 => X"96",  -- 150
        75796 => X"94",  -- 148
        75797 => X"81",  -- 129
        75798 => X"88",  -- 136
        75799 => X"89",  -- 137
        75800 => X"73",  -- 115
        75801 => X"67",  -- 103
        75802 => X"72",  -- 114
        75803 => X"6A",  -- 106
        75804 => X"58",  -- 88
        75805 => X"4D",  -- 77
        75806 => X"2C",  -- 44
        75807 => X"30",  -- 48
        75808 => X"21",  -- 33
        75809 => X"1D",  -- 29
        75810 => X"17",  -- 23
        75811 => X"15",  -- 21
        75812 => X"1B",  -- 27
        75813 => X"22",  -- 34
        75814 => X"25",  -- 37
        75815 => X"22",  -- 34
        75816 => X"2C",  -- 44
        75817 => X"18",  -- 24
        75818 => X"15",  -- 21
        75819 => X"30",  -- 48
        75820 => X"4F",  -- 79
        75821 => X"5C",  -- 92
        75822 => X"61",  -- 97
        75823 => X"65",  -- 101
        75824 => X"77",  -- 119
        75825 => X"78",  -- 120
        75826 => X"7E",  -- 126
        75827 => X"77",  -- 119
        75828 => X"6C",  -- 108
        75829 => X"6E",  -- 110
        75830 => X"76",  -- 118
        75831 => X"77",  -- 119
        75832 => X"61",  -- 97
        75833 => X"45",  -- 69
        75834 => X"44",  -- 68
        75835 => X"30",  -- 48
        75836 => X"33",  -- 51
        75837 => X"45",  -- 69
        75838 => X"4E",  -- 78
        75839 => X"83",  -- 131
        75840 => X"5E",  -- 94
        75841 => X"52",  -- 82
        75842 => X"4F",  -- 79
        75843 => X"53",  -- 83
        75844 => X"57",  -- 87
        75845 => X"60",  -- 96
        75846 => X"64",  -- 100
        75847 => X"5D",  -- 93
        75848 => X"48",  -- 72
        75849 => X"48",  -- 72
        75850 => X"44",  -- 68
        75851 => X"3C",  -- 60
        75852 => X"3F",  -- 63
        75853 => X"4D",  -- 77
        75854 => X"5A",  -- 90
        75855 => X"5F",  -- 95
        75856 => X"58",  -- 88
        75857 => X"5E",  -- 94
        75858 => X"5E",  -- 94
        75859 => X"5E",  -- 94
        75860 => X"61",  -- 97
        75861 => X"58",  -- 88
        75862 => X"4D",  -- 77
        75863 => X"4B",  -- 75
        75864 => X"50",  -- 80
        75865 => X"44",  -- 68
        75866 => X"51",  -- 81
        75867 => X"2B",  -- 43
        75868 => X"2F",  -- 47
        75869 => X"42",  -- 66
        75870 => X"52",  -- 82
        75871 => X"53",  -- 83
        75872 => X"59",  -- 89
        75873 => X"5F",  -- 95
        75874 => X"5E",  -- 94
        75875 => X"4D",  -- 77
        75876 => X"36",  -- 54
        75877 => X"2A",  -- 42
        75878 => X"2A",  -- 42
        75879 => X"2F",  -- 47
        75880 => X"44",  -- 68
        75881 => X"40",  -- 64
        75882 => X"44",  -- 68
        75883 => X"4B",  -- 75
        75884 => X"52",  -- 82
        75885 => X"4A",  -- 74
        75886 => X"43",  -- 67
        75887 => X"3B",  -- 59
        75888 => X"44",  -- 68
        75889 => X"4A",  -- 74
        75890 => X"51",  -- 81
        75891 => X"5E",  -- 94
        75892 => X"43",  -- 67
        75893 => X"38",  -- 56
        75894 => X"20",  -- 32
        75895 => X"2E",  -- 46
        75896 => X"23",  -- 35
        75897 => X"35",  -- 53
        75898 => X"2C",  -- 44
        75899 => X"13",  -- 19
        75900 => X"19",  -- 25
        75901 => X"33",  -- 51
        75902 => X"3E",  -- 62
        75903 => X"3B",  -- 59
        75904 => X"4C",  -- 76
        75905 => X"4A",  -- 74
        75906 => X"46",  -- 70
        75907 => X"47",  -- 71
        75908 => X"43",  -- 67
        75909 => X"30",  -- 48
        75910 => X"21",  -- 33
        75911 => X"27",  -- 39
        75912 => X"30",  -- 48
        75913 => X"37",  -- 55
        75914 => X"3F",  -- 63
        75915 => X"40",  -- 64
        75916 => X"3D",  -- 61
        75917 => X"38",  -- 56
        75918 => X"2E",  -- 46
        75919 => X"23",  -- 35
        75920 => X"1E",  -- 30
        75921 => X"30",  -- 48
        75922 => X"39",  -- 57
        75923 => X"31",  -- 49
        75924 => X"31",  -- 49
        75925 => X"39",  -- 57
        75926 => X"36",  -- 54
        75927 => X"29",  -- 41
        75928 => X"1F",  -- 31
        75929 => X"27",  -- 39
        75930 => X"29",  -- 41
        75931 => X"2E",  -- 46
        75932 => X"36",  -- 54
        75933 => X"2F",  -- 47
        75934 => X"22",  -- 34
        75935 => X"1F",  -- 31
        75936 => X"1D",  -- 29
        75937 => X"14",  -- 20
        75938 => X"17",  -- 23
        75939 => X"1F",  -- 31
        75940 => X"35",  -- 53
        75941 => X"3D",  -- 61
        75942 => X"30",  -- 48
        75943 => X"36",  -- 54
        75944 => X"34",  -- 52
        75945 => X"25",  -- 37
        75946 => X"2A",  -- 42
        75947 => X"2F",  -- 47
        75948 => X"21",  -- 33
        75949 => X"1F",  -- 31
        75950 => X"25",  -- 37
        75951 => X"20",  -- 32
        75952 => X"2F",  -- 47
        75953 => X"2D",  -- 45
        75954 => X"20",  -- 32
        75955 => X"1C",  -- 28
        75956 => X"29",  -- 41
        75957 => X"30",  -- 48
        75958 => X"2E",  -- 46
        75959 => X"2E",  -- 46
        75960 => X"32",  -- 50
        75961 => X"34",  -- 52
        75962 => X"37",  -- 55
        75963 => X"37",  -- 55
        75964 => X"34",  -- 52
        75965 => X"32",  -- 50
        75966 => X"33",  -- 51
        75967 => X"35",  -- 53
        75968 => X"3D",  -- 61
        75969 => X"3A",  -- 58
        75970 => X"37",  -- 55
        75971 => X"38",  -- 56
        75972 => X"3D",  -- 61
        75973 => X"42",  -- 66
        75974 => X"44",  -- 68
        75975 => X"43",  -- 67
        75976 => X"46",  -- 70
        75977 => X"42",  -- 66
        75978 => X"40",  -- 64
        75979 => X"40",  -- 64
        75980 => X"3B",  -- 59
        75981 => X"36",  -- 54
        75982 => X"37",  -- 55
        75983 => X"3D",  -- 61
        75984 => X"2E",  -- 46
        75985 => X"32",  -- 50
        75986 => X"38",  -- 56
        75987 => X"43",  -- 67
        75988 => X"41",  -- 65
        75989 => X"2B",  -- 43
        75990 => X"24",  -- 36
        75991 => X"33",  -- 51
        75992 => X"41",  -- 65
        75993 => X"38",  -- 56
        75994 => X"3D",  -- 61
        75995 => X"46",  -- 70
        75996 => X"42",  -- 66
        75997 => X"3D",  -- 61
        75998 => X"3D",  -- 61
        75999 => X"39",  -- 57
        76000 => X"39",  -- 57
        76001 => X"31",  -- 49
        76002 => X"36",  -- 54
        76003 => X"46",  -- 70
        76004 => X"48",  -- 72
        76005 => X"3B",  -- 59
        76006 => X"35",  -- 53
        76007 => X"3C",  -- 60
        76008 => X"34",  -- 52
        76009 => X"32",  -- 50
        76010 => X"39",  -- 57
        76011 => X"3F",  -- 63
        76012 => X"3F",  -- 63
        76013 => X"41",  -- 65
        76014 => X"44",  -- 68
        76015 => X"3C",  -- 60
        76016 => X"42",  -- 66
        76017 => X"4C",  -- 76
        76018 => X"50",  -- 80
        76019 => X"4E",  -- 78
        76020 => X"4E",  -- 78
        76021 => X"49",  -- 73
        76022 => X"44",  -- 68
        76023 => X"4B",  -- 75
        76024 => X"54",  -- 84
        76025 => X"55",  -- 85
        76026 => X"57",  -- 87
        76027 => X"58",  -- 88
        76028 => X"55",  -- 85
        76029 => X"46",  -- 70
        76030 => X"35",  -- 53
        76031 => X"29",  -- 41
        76032 => X"28",  -- 40
        76033 => X"36",  -- 54
        76034 => X"3F",  -- 63
        76035 => X"40",  -- 64
        76036 => X"44",  -- 68
        76037 => X"52",  -- 82
        76038 => X"63",  -- 99
        76039 => X"6B",  -- 107
        76040 => X"6A",  -- 106
        76041 => X"65",  -- 101
        76042 => X"5E",  -- 94
        76043 => X"59",  -- 89
        76044 => X"5B",  -- 91
        76045 => X"63",  -- 99
        76046 => X"6C",  -- 108
        76047 => X"73",  -- 115
        76048 => X"68",  -- 104
        76049 => X"59",  -- 89
        76050 => X"4B",  -- 75
        76051 => X"48",  -- 72
        76052 => X"50",  -- 80
        76053 => X"50",  -- 80
        76054 => X"42",  -- 66
        76055 => X"31",  -- 49
        76056 => X"39",  -- 57
        76057 => X"43",  -- 67
        76058 => X"40",  -- 64
        76059 => X"47",  -- 71
        76060 => X"4A",  -- 74
        76061 => X"3D",  -- 61
        76062 => X"40",  -- 64
        76063 => X"4A",  -- 74
        76064 => X"4C",  -- 76
        76065 => X"4C",  -- 76
        76066 => X"49",  -- 73
        76067 => X"47",  -- 71
        76068 => X"43",  -- 67
        76069 => X"43",  -- 67
        76070 => X"46",  -- 70
        76071 => X"48",  -- 72
        76072 => X"46",  -- 70
        76073 => X"4B",  -- 75
        76074 => X"4D",  -- 77
        76075 => X"46",  -- 70
        76076 => X"44",  -- 68
        76077 => X"49",  -- 73
        76078 => X"4B",  -- 75
        76079 => X"48",  -- 72
        76080 => X"3F",  -- 63
        76081 => X"45",  -- 69
        76082 => X"3F",  -- 63
        76083 => X"3C",  -- 60
        76084 => X"48",  -- 72
        76085 => X"50",  -- 80
        76086 => X"4E",  -- 78
        76087 => X"4D",  -- 77
        76088 => X"44",  -- 68
        76089 => X"48",  -- 72
        76090 => X"4F",  -- 79
        76091 => X"4B",  -- 75
        76092 => X"3C",  -- 60
        76093 => X"45",  -- 69
        76094 => X"43",  -- 67
        76095 => X"55",  -- 85
        76096 => X"7B",  -- 123
        76097 => X"55",  -- 85
        76098 => X"6D",  -- 109
        76099 => X"67",  -- 103
        76100 => X"59",  -- 89
        76101 => X"68",  -- 104
        76102 => X"58",  -- 88
        76103 => X"58",  -- 88
        76104 => X"5C",  -- 92
        76105 => X"4C",  -- 76
        76106 => X"5E",  -- 94
        76107 => X"47",  -- 71
        76108 => X"56",  -- 86
        76109 => X"2B",  -- 43
        76110 => X"34",  -- 52
        76111 => X"2D",  -- 45
        76112 => X"29",  -- 41
        76113 => X"4E",  -- 78
        76114 => X"5D",  -- 93
        76115 => X"6F",  -- 111
        76116 => X"80",  -- 128
        76117 => X"7F",  -- 127
        76118 => X"84",  -- 132
        76119 => X"63",  -- 99
        76120 => X"62",  -- 98
        76121 => X"63",  -- 99
        76122 => X"6C",  -- 108
        76123 => X"63",  -- 99
        76124 => X"51",  -- 81
        76125 => X"50",  -- 80
        76126 => X"32",  -- 50
        76127 => X"2F",  -- 47
        76128 => X"26",  -- 38
        76129 => X"2C",  -- 44
        76130 => X"2A",  -- 42
        76131 => X"23",  -- 35
        76132 => X"27",  -- 39
        76133 => X"40",  -- 64
        76134 => X"5C",  -- 92
        76135 => X"6B",  -- 107
        76136 => X"5F",  -- 95
        76137 => X"42",  -- 66
        76138 => X"3F",  -- 63
        76139 => X"60",  -- 96
        76140 => X"74",  -- 116
        76141 => X"6E",  -- 110
        76142 => X"76",  -- 118
        76143 => X"8F",  -- 143
        76144 => X"8D",  -- 141
        76145 => X"91",  -- 145
        76146 => X"93",  -- 147
        76147 => X"81",  -- 129
        76148 => X"66",  -- 102
        76149 => X"5E",  -- 94
        76150 => X"66",  -- 102
        76151 => X"69",  -- 105
        76152 => X"4A",  -- 74
        76153 => X"60",  -- 96
        76154 => X"85",  -- 133
        76155 => X"88",  -- 136
        76156 => X"91",  -- 145
        76157 => X"A0",  -- 160
        76158 => X"A0",  -- 160
        76159 => X"B8",  -- 184
        76160 => X"60",  -- 96
        76161 => X"53",  -- 83
        76162 => X"4D",  -- 77
        76163 => X"4E",  -- 78
        76164 => X"50",  -- 80
        76165 => X"5A",  -- 90
        76166 => X"63",  -- 99
        76167 => X"60",  -- 96
        76168 => X"62",  -- 98
        76169 => X"5E",  -- 94
        76170 => X"5B",  -- 91
        76171 => X"58",  -- 88
        76172 => X"5B",  -- 91
        76173 => X"60",  -- 96
        76174 => X"65",  -- 101
        76175 => X"68",  -- 104
        76176 => X"5B",  -- 91
        76177 => X"60",  -- 96
        76178 => X"5D",  -- 93
        76179 => X"56",  -- 86
        76180 => X"51",  -- 81
        76181 => X"43",  -- 67
        76182 => X"36",  -- 54
        76183 => X"35",  -- 53
        76184 => X"39",  -- 57
        76185 => X"36",  -- 54
        76186 => X"39",  -- 57
        76187 => X"2D",  -- 45
        76188 => X"32",  -- 50
        76189 => X"44",  -- 68
        76190 => X"51",  -- 81
        76191 => X"49",  -- 73
        76192 => X"4F",  -- 79
        76193 => X"57",  -- 87
        76194 => X"57",  -- 87
        76195 => X"46",  -- 70
        76196 => X"35",  -- 53
        76197 => X"31",  -- 49
        76198 => X"3A",  -- 58
        76199 => X"43",  -- 67
        76200 => X"56",  -- 86
        76201 => X"51",  -- 81
        76202 => X"55",  -- 85
        76203 => X"5C",  -- 92
        76204 => X"5A",  -- 90
        76205 => X"54",  -- 84
        76206 => X"4A",  -- 74
        76207 => X"40",  -- 64
        76208 => X"43",  -- 67
        76209 => X"4F",  -- 79
        76210 => X"48",  -- 72
        76211 => X"4E",  -- 78
        76212 => X"4A",  -- 74
        76213 => X"32",  -- 50
        76214 => X"23",  -- 35
        76215 => X"27",  -- 39
        76216 => X"2B",  -- 43
        76217 => X"3C",  -- 60
        76218 => X"36",  -- 54
        76219 => X"25",  -- 37
        76220 => X"31",  -- 49
        76221 => X"4B",  -- 75
        76222 => X"57",  -- 87
        76223 => X"57",  -- 87
        76224 => X"49",  -- 73
        76225 => X"4E",  -- 78
        76226 => X"49",  -- 73
        76227 => X"40",  -- 64
        76228 => X"36",  -- 54
        76229 => X"28",  -- 40
        76230 => X"22",  -- 34
        76231 => X"2D",  -- 45
        76232 => X"38",  -- 56
        76233 => X"3F",  -- 63
        76234 => X"47",  -- 71
        76235 => X"45",  -- 69
        76236 => X"41",  -- 65
        76237 => X"43",  -- 67
        76238 => X"3B",  -- 59
        76239 => X"2A",  -- 42
        76240 => X"1E",  -- 30
        76241 => X"23",  -- 35
        76242 => X"29",  -- 41
        76243 => X"2B",  -- 43
        76244 => X"2E",  -- 46
        76245 => X"33",  -- 51
        76246 => X"37",  -- 55
        76247 => X"38",  -- 56
        76248 => X"35",  -- 53
        76249 => X"39",  -- 57
        76250 => X"32",  -- 50
        76251 => X"2D",  -- 45
        76252 => X"37",  -- 55
        76253 => X"3C",  -- 60
        76254 => X"33",  -- 51
        76255 => X"2D",  -- 45
        76256 => X"31",  -- 49
        76257 => X"1C",  -- 28
        76258 => X"15",  -- 21
        76259 => X"1E",  -- 30
        76260 => X"3C",  -- 60
        76261 => X"46",  -- 70
        76262 => X"30",  -- 48
        76263 => X"2C",  -- 44
        76264 => X"32",  -- 50
        76265 => X"25",  -- 37
        76266 => X"2B",  -- 43
        76267 => X"2C",  -- 44
        76268 => X"1C",  -- 28
        76269 => X"23",  -- 35
        76270 => X"32",  -- 50
        76271 => X"2C",  -- 44
        76272 => X"2F",  -- 47
        76273 => X"31",  -- 49
        76274 => X"27",  -- 39
        76275 => X"21",  -- 33
        76276 => X"2A",  -- 42
        76277 => X"33",  -- 51
        76278 => X"36",  -- 54
        76279 => X"3B",  -- 59
        76280 => X"39",  -- 57
        76281 => X"3C",  -- 60
        76282 => X"3E",  -- 62
        76283 => X"3C",  -- 60
        76284 => X"3A",  -- 58
        76285 => X"39",  -- 57
        76286 => X"3A",  -- 58
        76287 => X"3B",  -- 59
        76288 => X"37",  -- 55
        76289 => X"37",  -- 55
        76290 => X"3A",  -- 58
        76291 => X"3E",  -- 62
        76292 => X"46",  -- 70
        76293 => X"4A",  -- 74
        76294 => X"4A",  -- 74
        76295 => X"49",  -- 73
        76296 => X"4A",  -- 74
        76297 => X"41",  -- 65
        76298 => X"3D",  -- 61
        76299 => X"40",  -- 64
        76300 => X"3F",  -- 63
        76301 => X"38",  -- 56
        76302 => X"35",  -- 53
        76303 => X"38",  -- 56
        76304 => X"37",  -- 55
        76305 => X"42",  -- 66
        76306 => X"43",  -- 67
        76307 => X"44",  -- 68
        76308 => X"47",  -- 71
        76309 => X"3D",  -- 61
        76310 => X"36",  -- 54
        76311 => X"3F",  -- 63
        76312 => X"36",  -- 54
        76313 => X"32",  -- 50
        76314 => X"3C",  -- 60
        76315 => X"45",  -- 69
        76316 => X"40",  -- 64
        76317 => X"43",  -- 67
        76318 => X"45",  -- 69
        76319 => X"3A",  -- 58
        76320 => X"3D",  -- 61
        76321 => X"38",  -- 56
        76322 => X"3F",  -- 63
        76323 => X"4C",  -- 76
        76324 => X"4B",  -- 75
        76325 => X"3B",  -- 59
        76326 => X"33",  -- 51
        76327 => X"35",  -- 53
        76328 => X"37",  -- 55
        76329 => X"39",  -- 57
        76330 => X"42",  -- 66
        76331 => X"45",  -- 69
        76332 => X"40",  -- 64
        76333 => X"41",  -- 65
        76334 => X"49",  -- 73
        76335 => X"49",  -- 73
        76336 => X"4A",  -- 74
        76337 => X"51",  -- 81
        76338 => X"4F",  -- 79
        76339 => X"4B",  -- 75
        76340 => X"4E",  -- 78
        76341 => X"4C",  -- 76
        76342 => X"4A",  -- 74
        76343 => X"51",  -- 81
        76344 => X"41",  -- 65
        76345 => X"4F",  -- 79
        76346 => X"57",  -- 87
        76347 => X"51",  -- 81
        76348 => X"45",  -- 69
        76349 => X"3D",  -- 61
        76350 => X"34",  -- 52
        76351 => X"2C",  -- 44
        76352 => X"31",  -- 49
        76353 => X"3B",  -- 59
        76354 => X"42",  -- 66
        76355 => X"41",  -- 65
        76356 => X"47",  -- 71
        76357 => X"55",  -- 85
        76358 => X"62",  -- 98
        76359 => X"66",  -- 102
        76360 => X"61",  -- 97
        76361 => X"5D",  -- 93
        76362 => X"58",  -- 88
        76363 => X"54",  -- 84
        76364 => X"54",  -- 84
        76365 => X"5F",  -- 95
        76366 => X"6D",  -- 109
        76367 => X"78",  -- 120
        76368 => X"70",  -- 112
        76369 => X"61",  -- 97
        76370 => X"54",  -- 84
        76371 => X"52",  -- 82
        76372 => X"5A",  -- 90
        76373 => X"5D",  -- 93
        76374 => X"5B",  -- 91
        76375 => X"57",  -- 87
        76376 => X"50",  -- 80
        76377 => X"47",  -- 71
        76378 => X"42",  -- 66
        76379 => X"48",  -- 72
        76380 => X"57",  -- 87
        76381 => X"50",  -- 80
        76382 => X"42",  -- 66
        76383 => X"53",  -- 83
        76384 => X"50",  -- 80
        76385 => X"4F",  -- 79
        76386 => X"4B",  -- 75
        76387 => X"49",  -- 73
        76388 => X"47",  -- 71
        76389 => X"48",  -- 72
        76390 => X"49",  -- 73
        76391 => X"4B",  -- 75
        76392 => X"4B",  -- 75
        76393 => X"48",  -- 72
        76394 => X"4C",  -- 76
        76395 => X"54",  -- 84
        76396 => X"53",  -- 83
        76397 => X"4B",  -- 75
        76398 => X"4A",  -- 74
        76399 => X"50",  -- 80
        76400 => X"45",  -- 69
        76401 => X"51",  -- 81
        76402 => X"4E",  -- 78
        76403 => X"47",  -- 71
        76404 => X"4A",  -- 74
        76405 => X"49",  -- 73
        76406 => X"41",  -- 65
        76407 => X"3D",  -- 61
        76408 => X"3D",  -- 61
        76409 => X"4F",  -- 79
        76410 => X"54",  -- 84
        76411 => X"45",  -- 69
        76412 => X"35",  -- 53
        76413 => X"4D",  -- 77
        76414 => X"45",  -- 69
        76415 => X"45",  -- 69
        76416 => X"60",  -- 96
        76417 => X"54",  -- 84
        76418 => X"5D",  -- 93
        76419 => X"51",  -- 81
        76420 => X"4A",  -- 74
        76421 => X"52",  -- 82
        76422 => X"45",  -- 69
        76423 => X"48",  -- 72
        76424 => X"5B",  -- 91
        76425 => X"4C",  -- 76
        76426 => X"59",  -- 89
        76427 => X"3F",  -- 63
        76428 => X"59",  -- 89
        76429 => X"2E",  -- 46
        76430 => X"35",  -- 53
        76431 => X"29",  -- 41
        76432 => X"3E",  -- 62
        76433 => X"56",  -- 86
        76434 => X"58",  -- 88
        76435 => X"58",  -- 88
        76436 => X"72",  -- 114
        76437 => X"6A",  -- 106
        76438 => X"75",  -- 117
        76439 => X"47",  -- 71
        76440 => X"5C",  -- 92
        76441 => X"63",  -- 99
        76442 => X"61",  -- 97
        76443 => X"60",  -- 96
        76444 => X"4F",  -- 79
        76445 => X"59",  -- 89
        76446 => X"4C",  -- 76
        76447 => X"4E",  -- 78
        76448 => X"51",  -- 81
        76449 => X"49",  -- 73
        76450 => X"45",  -- 69
        76451 => X"52",  -- 82
        76452 => X"6A",  -- 106
        76453 => X"81",  -- 129
        76454 => X"85",  -- 133
        76455 => X"7F",  -- 127
        76456 => X"76",  -- 118
        76457 => X"68",  -- 104
        76458 => X"68",  -- 104
        76459 => X"79",  -- 121
        76460 => X"82",  -- 130
        76461 => X"7F",  -- 127
        76462 => X"87",  -- 135
        76463 => X"99",  -- 153
        76464 => X"9A",  -- 154
        76465 => X"8B",  -- 139
        76466 => X"7B",  -- 123
        76467 => X"68",  -- 104
        76468 => X"5C",  -- 92
        76469 => X"67",  -- 103
        76470 => X"7A",  -- 122
        76471 => X"80",  -- 128
        76472 => X"8A",  -- 138
        76473 => X"AF",  -- 175
        76474 => X"BA",  -- 186
        76475 => X"A4",  -- 164
        76476 => X"A0",  -- 160
        76477 => X"A7",  -- 167
        76478 => X"98",  -- 152
        76479 => X"82",  -- 130
        76480 => X"7A",  -- 122
        76481 => X"6D",  -- 109
        76482 => X"67",  -- 103
        76483 => X"66",  -- 102
        76484 => X"65",  -- 101
        76485 => X"6D",  -- 109
        76486 => X"74",  -- 116
        76487 => X"70",  -- 112
        76488 => X"65",  -- 101
        76489 => X"63",  -- 99
        76490 => X"67",  -- 103
        76491 => X"6D",  -- 109
        76492 => X"71",  -- 113
        76493 => X"6F",  -- 111
        76494 => X"6A",  -- 106
        76495 => X"67",  -- 103
        76496 => X"6B",  -- 107
        76497 => X"6F",  -- 111
        76498 => X"65",  -- 101
        76499 => X"58",  -- 88
        76500 => X"52",  -- 82
        76501 => X"48",  -- 72
        76502 => X"42",  -- 66
        76503 => X"48",  -- 72
        76504 => X"42",  -- 66
        76505 => X"44",  -- 68
        76506 => X"40",  -- 64
        76507 => X"49",  -- 73
        76508 => X"51",  -- 81
        76509 => X"64",  -- 100
        76510 => X"6F",  -- 111
        76511 => X"61",  -- 97
        76512 => X"58",  -- 88
        76513 => X"65",  -- 101
        76514 => X"66",  -- 102
        76515 => X"54",  -- 84
        76516 => X"41",  -- 65
        76517 => X"41",  -- 65
        76518 => X"52",  -- 82
        76519 => X"60",  -- 96
        76520 => X"5F",  -- 95
        76521 => X"59",  -- 89
        76522 => X"5C",  -- 92
        76523 => X"66",  -- 102
        76524 => X"64",  -- 100
        76525 => X"66",  -- 102
        76526 => X"62",  -- 98
        76527 => X"5A",  -- 90
        76528 => X"5A",  -- 90
        76529 => X"61",  -- 97
        76530 => X"4D",  -- 77
        76531 => X"48",  -- 72
        76532 => X"65",  -- 101
        76533 => X"47",  -- 71
        76534 => X"3D",  -- 61
        76535 => X"2A",  -- 42
        76536 => X"3A",  -- 58
        76537 => X"44",  -- 68
        76538 => X"3E",  -- 62
        76539 => X"35",  -- 53
        76540 => X"42",  -- 66
        76541 => X"56",  -- 86
        76542 => X"5F",  -- 95
        76543 => X"61",  -- 97
        76544 => X"5A",  -- 90
        76545 => X"64",  -- 100
        76546 => X"5F",  -- 95
        76547 => X"4F",  -- 79
        76548 => X"40",  -- 64
        76549 => X"35",  -- 53
        76550 => X"38",  -- 56
        76551 => X"47",  -- 71
        76552 => X"49",  -- 73
        76553 => X"4E",  -- 78
        76554 => X"53",  -- 83
        76555 => X"4C",  -- 76
        76556 => X"48",  -- 72
        76557 => X"4F",  -- 79
        76558 => X"49",  -- 73
        76559 => X"32",  -- 50
        76560 => X"34",  -- 52
        76561 => X"2E",  -- 46
        76562 => X"31",  -- 49
        76563 => X"3E",  -- 62
        76564 => X"45",  -- 69
        76565 => X"45",  -- 69
        76566 => X"4F",  -- 79
        76567 => X"5E",  -- 94
        76568 => X"54",  -- 84
        76569 => X"52",  -- 82
        76570 => X"3F",  -- 63
        76571 => X"32",  -- 50
        76572 => X"3F",  -- 63
        76573 => X"4D",  -- 77
        76574 => X"49",  -- 73
        76575 => X"40",  -- 64
        76576 => X"3A",  -- 58
        76577 => X"34",  -- 52
        76578 => X"32",  -- 50
        76579 => X"2B",  -- 43
        76580 => X"34",  -- 52
        76581 => X"3B",  -- 59
        76582 => X"33",  -- 51
        76583 => X"3C",  -- 60
        76584 => X"37",  -- 55
        76585 => X"2C",  -- 44
        76586 => X"36",  -- 54
        76587 => X"37",  -- 55
        76588 => X"28",  -- 40
        76589 => X"34",  -- 52
        76590 => X"45",  -- 69
        76591 => X"3B",  -- 59
        76592 => X"39",  -- 57
        76593 => X"3F",  -- 63
        76594 => X"37",  -- 55
        76595 => X"2E",  -- 46
        76596 => X"32",  -- 50
        76597 => X"3C",  -- 60
        76598 => X"44",  -- 68
        76599 => X"4E",  -- 78
        76600 => X"44",  -- 68
        76601 => X"47",  -- 71
        76602 => X"49",  -- 73
        76603 => X"48",  -- 72
        76604 => X"46",  -- 70
        76605 => X"47",  -- 71
        76606 => X"4A",  -- 74
        76607 => X"4B",  -- 75
        76608 => X"41",  -- 65
        76609 => X"44",  -- 68
        76610 => X"48",  -- 72
        76611 => X"4E",  -- 78
        76612 => X"52",  -- 82
        76613 => X"54",  -- 84
        76614 => X"4F",  -- 79
        76615 => X"4B",  -- 75
        76616 => X"4E",  -- 78
        76617 => X"43",  -- 67
        76618 => X"40",  -- 64
        76619 => X"4A",  -- 74
        76620 => X"53",  -- 83
        76621 => X"51",  -- 81
        76622 => X"4E",  -- 78
        76623 => X"50",  -- 80
        76624 => X"4A",  -- 74
        76625 => X"59",  -- 89
        76626 => X"4F",  -- 79
        76627 => X"43",  -- 67
        76628 => X"4C",  -- 76
        76629 => X"52",  -- 82
        76630 => X"4F",  -- 79
        76631 => X"53",  -- 83
        76632 => X"4B",  -- 75
        76633 => X"49",  -- 73
        76634 => X"50",  -- 80
        76635 => X"4A",  -- 74
        76636 => X"39",  -- 57
        76637 => X"40",  -- 64
        76638 => X"54",  -- 84
        76639 => X"54",  -- 84
        76640 => X"4F",  -- 79
        76641 => X"4D",  -- 77
        76642 => X"55",  -- 85
        76643 => X"5E",  -- 94
        76644 => X"59",  -- 89
        76645 => X"48",  -- 72
        76646 => X"3D",  -- 61
        76647 => X"3D",  -- 61
        76648 => X"4C",  -- 76
        76649 => X"40",  -- 64
        76650 => X"40",  -- 64
        76651 => X"49",  -- 73
        76652 => X"50",  -- 80
        76653 => X"59",  -- 89
        76654 => X"5C",  -- 92
        76655 => X"55",  -- 85
        76656 => X"58",  -- 88
        76657 => X"5C",  -- 92
        76658 => X"55",  -- 85
        76659 => X"4F",  -- 79
        76660 => X"52",  -- 82
        76661 => X"50",  -- 80
        76662 => X"51",  -- 81
        76663 => X"59",  -- 89
        76664 => X"58",  -- 88
        76665 => X"55",  -- 85
        76666 => X"54",  -- 84
        76667 => X"57",  -- 87
        76668 => X"5A",  -- 90
        76669 => X"5B",  -- 91
        76670 => X"5A",  -- 90
        76671 => X"57",  -- 87
        76672 => X"49",  -- 73
        76673 => X"4D",  -- 77
        76674 => X"4D",  -- 77
        76675 => X"49",  -- 73
        76676 => X"51",  -- 81
        76677 => X"5F",  -- 95
        76678 => X"66",  -- 102
        76679 => X"65",  -- 101
        76680 => X"6A",  -- 106
        76681 => X"68",  -- 104
        76682 => X"63",  -- 99
        76683 => X"5F",  -- 95
        76684 => X"5F",  -- 95
        76685 => X"6C",  -- 108
        76686 => X"7E",  -- 126
        76687 => X"8B",  -- 139
        76688 => X"84",  -- 132
        76689 => X"74",  -- 116
        76690 => X"62",  -- 98
        76691 => X"5F",  -- 95
        76692 => X"63",  -- 99
        76693 => X"63",  -- 99
        76694 => X"67",  -- 103
        76695 => X"6C",  -- 108
        76696 => X"51",  -- 81
        76697 => X"48",  -- 72
        76698 => X"50",  -- 80
        76699 => X"4F",  -- 79
        76700 => X"55",  -- 85
        76701 => X"4C",  -- 76
        76702 => X"3F",  -- 63
        76703 => X"63",  -- 99
        76704 => X"5D",  -- 93
        76705 => X"5C",  -- 92
        76706 => X"57",  -- 87
        76707 => X"54",  -- 84
        76708 => X"51",  -- 81
        76709 => X"51",  -- 81
        76710 => X"51",  -- 81
        76711 => X"52",  -- 82
        76712 => X"53",  -- 83
        76713 => X"3F",  -- 63
        76714 => X"42",  -- 66
        76715 => X"5C",  -- 92
        76716 => X"67",  -- 103
        76717 => X"57",  -- 87
        76718 => X"4D",  -- 77
        76719 => X"54",  -- 84
        76720 => X"54",  -- 84
        76721 => X"60",  -- 96
        76722 => X"5B",  -- 91
        76723 => X"4F",  -- 79
        76724 => X"4F",  -- 79
        76725 => X"52",  -- 82
        76726 => X"53",  -- 83
        76727 => X"57",  -- 87
        76728 => X"5A",  -- 90
        76729 => X"50",  -- 80
        76730 => X"52",  -- 82
        76731 => X"61",  -- 97
        76732 => X"52",  -- 82
        76733 => X"50",  -- 80
        76734 => X"40",  -- 64
        76735 => X"55",  -- 85
        76736 => X"56",  -- 86
        76737 => X"6E",  -- 110
        76738 => X"65",  -- 101
        76739 => X"55",  -- 85
        76740 => X"59",  -- 89
        76741 => X"56",  -- 86
        76742 => X"51",  -- 81
        76743 => X"56",  -- 86
        76744 => X"6B",  -- 107
        76745 => X"62",  -- 98
        76746 => X"5A",  -- 90
        76747 => X"50",  -- 80
        76748 => X"5E",  -- 94
        76749 => X"52",  -- 82
        76750 => X"4B",  -- 75
        76751 => X"43",  -- 67
        76752 => X"4F",  -- 79
        76753 => X"68",  -- 104
        76754 => X"75",  -- 117
        76755 => X"70",  -- 112
        76756 => X"7B",  -- 123
        76757 => X"60",  -- 96
        76758 => X"8B",  -- 139
        76759 => X"81",  -- 129
        76760 => X"72",  -- 114
        76761 => X"76",  -- 118
        76762 => X"68",  -- 104
        76763 => X"6C",  -- 108
        76764 => X"5D",  -- 93
        76765 => X"6C",  -- 108
        76766 => X"71",  -- 113
        76767 => X"7D",  -- 125
        76768 => X"6E",  -- 110
        76769 => X"70",  -- 112
        76770 => X"7D",  -- 125
        76771 => X"8F",  -- 143
        76772 => X"99",  -- 153
        76773 => X"9A",  -- 154
        76774 => X"9A",  -- 154
        76775 => X"9E",  -- 158
        76776 => X"8D",  -- 141
        76777 => X"8B",  -- 139
        76778 => X"86",  -- 134
        76779 => X"8B",  -- 139
        76780 => X"A1",  -- 161
        76781 => X"AE",  -- 174
        76782 => X"99",  -- 153
        76783 => X"76",  -- 118
        76784 => X"88",  -- 136
        76785 => X"89",  -- 137
        76786 => X"92",  -- 146
        76787 => X"97",  -- 151
        76788 => X"9C",  -- 156
        76789 => X"AD",  -- 173
        76790 => X"BD",  -- 189
        76791 => X"BF",  -- 191
        76792 => X"A5",  -- 165
        76793 => X"BC",  -- 188
        76794 => X"B5",  -- 181
        76795 => X"A2",  -- 162
        76796 => X"96",  -- 150
        76797 => X"8F",  -- 143
        76798 => X"97",  -- 151
        76799 => X"99"   -- 153
    );
    
begin
    
    process(clk)
    begin
        if rising_edge(clk) then
            if re = '1' then
                dout_reg <= mem(to_integer(unsigned(addr)));
            end if;
        end if;
    end process;

    -- Output assignment
    dout <= dout_reg;
    
end architecture rtl;
